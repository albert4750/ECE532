localparam bit signed [0:146][7:0] Input4 = '{27, 103, -101, -99, -2, -56, -53, -31, 78, -90, -117, 74, 118, -39, -96, 50, -88, 70, -98, 22, -5, -53, -93, 84, 68, -65, -124, 49, -12, 29, 63, -67, -37, -17, 83, -24, -38, -102, -55, 50, 95, -34, -111, 71, -72, 115, -93, 73, 92, -81, -80, -9, 71, -11, -61, -5, 71, -66, 72, -91, -123, -31, -73, 92, 46, -90, -79, -120, -6, 65, -62, -66, -112, 61, 66, -117, 31, 10, -108, -28, -114, -8, -76, 71, 29, 5, -114, -14, 110, 79, -77, -96, 23, 121, -37, -122, 73, -8, -63, -53, -41, 124, 70, -88, 60, -92, 12, 35, -66, 69, -66, 58, -52, -110, 0, -127, 84, 77, -38, -16, -21, 21, -50, -115, 104, -61, -23, 17, -123, -102, 63, 27, 107, 109, 41, -115, -83, 48, -72, -70, -111, 86, -33, 89, 92, 77, 7};
