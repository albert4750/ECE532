localparam bit signed [0:15][7:0] Output3 = '{32, -127, -120, -53, 95, 101, -113, -127, 126, -47, 16, 6, 14, 71, -48, -1};
