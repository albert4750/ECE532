localparam bit signed [0:2][0:7][0:2][0:2][24:0] Weight3 = '{
    '{'{'{-25'd155543, 25'd224477, -25'd174986}, '{25'd28281, 25'd113122, 25'd0}, '{-25'd81307, 25'd51259, 25'd15908}}, '{'{-25'd21210, 25'd19443, -25'd76004}, '{-25'd91912, -25'd104285, 25'd10605}, '{25'd21210, 25'd31816, -25'd79539}}, '{'{-25'd17675, 25'd91912, 25'd68934}, '{25'd125495, 25'd54794, 25'd144938}, '{25'd106052, 25'd44188, 25'd42421}}, '{'{25'd125495, -25'd70701, -25'd90144}, '{-25'd144938, -25'd70701, -25'd26513}, '{-25'd40653, -25'd10605, -25'd45956}}, '{'{25'd97215, 25'd106052, 25'd21210}, '{25'd83074, 25'd1768, 25'd45956}, '{25'd61864, -25'd22978, -25'd30048}}, '{'{25'd47724, 25'd37118, -25'd37118}, '{-25'd21210, -25'd35351, 25'd35351}, '{-25'd49491, -25'd67166, 25'd30048}}, '{'{-25'd49491, -25'd60096, -25'd84842}, '{25'd14140, 25'd7070, -25'd44188}, '{25'd74237, 25'd81307, -25'd1768}}, '{'{-25'd37118, 25'd47724, 25'd84842}, '{25'd136100, 25'd53026, -25'd35351}, '{25'd7070, 25'd113122, -25'd1768}}},
    '{'{'{-25'd205474, 25'd207783, -25'd64644}, '{25'd293204, 25'd106200, 25'd2309}, '{-25'd161609, 25'd6926, -25'd85422}}, '{'{-25'd83113, -25'd87730, 25'd53100}, '{-25'd60026, -25'd62335, 25'd20778}, '{-25'd36939, 25'd27704, 25'd23087}}, '{'{-25'd46174, 25'd73878, -25'd25396}, '{-25'd64644, -25'd25396, 25'd18470}, '{25'd66952, 25'd106200, -25'd80804}}, '{'{25'd145448, 25'd50791, -25'd55409}, '{-25'd30013, -25'd32322, 25'd233178}, '{-25'd6926, -25'd66952, 25'd101583}}, '{'{25'd27704, -25'd2309, 25'd96965}, '{-25'd39248, -25'd30013, 25'd39248}, '{25'd73878, 25'd73878, -25'd6926}}, '{'{-25'd57717, 25'd110817, 25'd133904}, '{25'd55409, 25'd55409, 25'd53100}, '{-25'd62335, 25'd9235, 25'd217017}}, '{'{-25'd32322, -25'd80804, -25'd73878}, '{25'd41557, 25'd69261, 25'd76187}, '{25'd23087, -25'd13852, 25'd2309}}, '{'{-25'd13852, 25'd30013, 25'd133904}, '{25'd9235, -25'd39248, -25'd36939}, '{-25'd25396, 25'd87730, 25'd39248}}},
    '{'{'{-25'd125534, 25'd20542, -25'd141511}, '{-25'd269327, -25'd52496, -25'd100427}, '{-25'd223678, 25'd289869, -25'd205419}}, '{'{-25'd36519, -25'd20542, -25'd130099}, '{-25'd6847, -25'd102709, -25'd114121}, '{-25'd155205, -25'd9130, -25'd104992}}, '{'{25'd111839, 25'd18259, 25'd6847}, '{25'd114121, 25'd219113, 25'd102709}, '{-25'd11412, 25'd120969, -25'd9130}}, '{'{25'd15977, 25'd31954, 25'd15977}, '{25'd155205, 25'd66190, 25'd95862}, '{-25'd102709, 25'd13695, 25'd11412}}, '{'{-25'd43366, -25'd15977, 25'd11412}, '{25'd114121, 25'd95862, 25'd123251}, '{25'd127816, 25'd22824, 25'd45649}}, '{'{-25'd34236, -25'd70755, -25'd66190}, '{-25'd89015, -25'd98144, 25'd4565}, '{-25'd109557, 25'd29672, -25'd70755}}, '{'{-25'd2282, 25'd54778, -25'd79885}, '{-25'd38801, -25'd52496, -25'd38801}, '{25'd45649, -25'd2282, -25'd2282}}, '{'{25'd114121, 25'd15977, 25'd31954}, '{25'd38801, -25'd25107, 25'd100427}, '{-25'd27389, 25'd6847, 25'd98144}}}
};
