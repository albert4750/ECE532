localparam bit signed [0:2][0:26][19:0] Input5 = '{
    '{-20'd45, 20'd49, -20'd87, -20'd35, 20'd46, 20'd21, 20'd73, -20'd39, 20'd114, 20'd96, 20'd91, -20'd55, -20'd100, 20'd107, 20'd81, -20'd23, 20'd58, 20'd0, 20'd86, -20'd65, -20'd112, -20'd22, 20'd36, -20'd34, -20'd104, -20'd12, 20'd63},
    '{20'd67, -20'd77, 20'd8, 20'd56, -20'd37, -20'd35, -20'd5, 20'd110, -20'd41, 20'd32, 20'd19, -20'd56, 20'd71, -20'd41, -20'd115, -20'd70, -20'd47, -20'd8, -20'd12, 20'd55, -20'd64, 20'd75, 20'd92, 20'd36, -20'd103, -20'd96, 20'd42},
    '{-20'd114, 20'd86, -20'd100, -20'd108, 20'd82, -20'd60, -20'd106, 20'd99, -20'd6, -20'd45, 20'd7, 20'd72, -20'd67, 20'd13, -20'd123, -20'd128, 20'd8, 20'd79, 20'd79, 20'd53, 20'd11, -20'd124, 20'd39, -20'd36, 20'd45, -20'd102, -20'd54}
};
