localparam bit signed [0:26][19:0] Output8 = '{20'd87, -20'd139, 20'd140, 20'd179, 20'd204, 20'd9, 20'd66, -20'd173, -20'd47, -20'd51, 20'd93, 20'd43, 20'd66, 20'd82, 20'd152, 20'd116, -20'd40, -20'd49, -20'd112, -20'd28, -20'd131, 20'd63, 20'd23, 20'd27, 20'd79, -20'd20, 20'd76};
