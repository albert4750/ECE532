localparam bit signed [0:7][0:2][0:2][0:2][24:0] Weight1 = '{
    '{'{'{25'd1214, -25'd1581, 25'd1166}, '{25'd256, 25'd958, 25'd830}, '{25'd2028, -25'd591, 25'd48}}, '{'{25'd447, 25'd1549, 25'd319}, '{-25'd240, -25'd1517, -25'd240}, '{-25'd287, -25'd272, -25'd735}}, '{'{25'd1613, 25'd974, -25'd830}, '{25'd1086, -25'd495, -25'd591}, '{25'd112, 25'd0, 25'd687}}},
    '{'{'{25'd452, -25'd291, -25'd2067}, '{25'd0, -25'd1243, 25'd1825}, '{25'd1308, 25'd452, -25'd711}}, '{'{25'd81, -25'd323, 25'd775}, '{-25'd581, -25'd1050, -25'd646}, '{-25'd226, 25'd1114, -25'd824}}, '{'{25'd65, -25'd791, -25'd1470}, '{-25'd1308, -25'd16, -25'd630}, '{-25'd549, -25'd872, 25'd194}}},
    '{'{'{25'd1311, 25'd1677, -25'd1053}, '{25'd258, 25'd1612, -25'd21}, '{25'd838, -25'd881, -25'd473}}, '{'{25'd1763, -25'd2085, 25'd709}, '{25'd2537, 25'd2666, 25'd473}, '{-25'd473, 25'd1741, -25'd86}}, '{'{25'd817, 25'd473, -25'd1096}, '{25'd1397, -25'd666, -25'd236}, '{-25'd1935, -25'd2730, -25'd451}}},
    '{'{'{-25'd306, -25'd274, -25'd1368}, '{25'd998, 25'd1594, 25'd1755}, '{-25'd2061, 25'd258, -25'd1900}}, '{'{-25'd757, 25'd419, -25'd2061}, '{25'd1497, 25'd1417, -25'd177}, '{-25'd1481, 25'd1755, -25'd2029}}, '{'{-25'd1594, 25'd547, -25'd16}, '{25'd402, 25'd1771, 25'd837}, '{25'd563, -25'd724, -25'd1014}}},
    '{'{'{-25'd469, -25'd566, -25'd1585}, '{25'd1132, -25'd1342, -25'd16}, '{-25'd1035, -25'd356, 25'd356}}, '{'{25'd744, -25'd1504, 25'd663}, '{-25'd1650, -25'd696, 25'd809}, '{25'd615, 25'd566, -25'd2070}}, '{'{25'd712, 25'd485, 25'd582}, '{-25'd906, -25'd1520, -25'd1747}, '{-25'd1375, 25'd809, 25'd598}}},
    '{'{'{-25'd1407, -25'd1139, 25'd1306}, '{-25'd100, 25'd1407, 25'd268}, '{25'd234, 25'd1675, 25'd268}}, '{'{-25'd4287, -25'd100, 25'd804}, '{-25'd3517, -25'd67, -25'd703}, '{-25'd1139, 25'd1407, -25'd1541}}, '{'{-25'd1708, 25'd2110, -25'd1574}, '{-25'd3082, -25'd670, -25'd1708}, '{-25'd703, 25'd2311, 25'd100}}},
    '{'{'{25'd445, 25'd801, -25'd1038}, '{25'd2136, 25'd2432, 25'd2314}, '{25'd3767, 25'd1187, -25'd623}}, '{'{25'd1127, -25'd534, -25'd267}, '{-25'd59, 25'd1928, 25'd2077}, '{-25'd1246, 25'd1602, -25'd1424}}, '{'{25'd2047, 25'd0, -25'd534}, '{-25'd237, 25'd415, -25'd1276}, '{-25'd801, 25'd1543, -25'd890}}},
    '{'{'{25'd200, 25'd89, -25'd1469}, '{25'd1202, -25'd801, 25'd423}, '{-25'd534, -25'd668, -25'd801}}, '{'{25'd267, 25'd2115, 25'd757}, '{25'd2382, 25'd868, -25'd245}, '{25'd1202, 25'd1358, 25'd1046}}, '{'{-25'd1135, 25'd423, -25'd1135}, '{-25'd89, 25'd2827, 25'd2048}, '{25'd690, 25'd1736, -25'd668}}}
};
