localparam bit signed [0:26][19:0] Output0 = '{-20'd60, -20'd228, -20'd164, 20'd19, 20'd75, 20'd133, 20'd182, 20'd216, 20'd25, 20'd195, -20'd101, 20'd61, -20'd122, -20'd87, -20'd87, 20'd212, -20'd66, 20'd132, -20'd259, 20'd188, 20'd237, -20'd186, -20'd51, -20'd46, 20'd2, -20'd252, 20'd152};
