localparam bit signed [0:31][47:0] Bias2 = '{48'd26381, -48'd76462, -48'd38935, -48'd49971, -48'd91487, -48'd49720, 48'd16850, 48'd38609, -48'd41667, -48'd37669, 48'd23914, -48'd6143, 48'd104319, 48'd87573, 48'd80509, -48'd126796, 48'd44692, -48'd67259, 48'd60468, 48'd42414, 48'd115279, -48'd85135, 48'd307048, 48'd121567, -48'd62958, -48'd146434, 48'd70640, 48'd91461, -48'd4797, 48'd12983, -48'd41440, 48'd28064};
