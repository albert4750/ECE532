localparam bit signed [0:46][15:0] Input2 = '{-16'd13428, -16'd25372, 16'd3898, 16'd20353, -16'd18063, 16'd23680, -16'd11481, 16'd29720, -16'd7494, -16'd16092, -16'd1693, 16'd25413, 16'd14470, 16'd20483, -16'd27422, -16'd9351, 16'd4776, -16'd1604, -16'd19039, -16'd8932, 16'd23364, -16'd28646, -16'd32032, -16'd5896, 16'd4461, -16'd14413, -16'd21303, -16'd19019, 16'd8389, 16'd13217, 16'd1671, 16'd27261, 16'd606, -16'd14264, 16'd12534, 16'd23380, 16'd25735, 16'd18115, 16'd26837, -16'd16933, -16'd24980, 16'd19779, 16'd6246, -16'd8364, -16'd5817, -16'd7597, 16'd5343};
