localparam bit signed [0:26][19:0] Output9 = '{-20'd59, 20'd66, 20'd95, 20'd4, 20'd38, 20'd44, -20'd20, -20'd243, 20'd191, 20'd148, -20'd26, 20'd64, -20'd156, 20'd233, -20'd117, 20'd122, -20'd111, -20'd53, 20'd84, 20'd282, 20'd54, -20'd122, 20'd120, 20'd43, 20'd123, 20'd177, 20'd49};
