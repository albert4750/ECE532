localparam bit signed [0:15][7:0] Output2 = '{-35, -21, -104, 32, -111, 61, -103, 40, 113, 29, -32, 20, -110, -11, 54, -108};
