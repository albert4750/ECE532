localparam bit signed [0:2][47:0] Bias3 = '{48'd1388, 48'd1341, 48'd1386};
