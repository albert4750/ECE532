localparam bit signed [0:15][7:0] Output0 = '{14, 92, 34, 5, 113, 14, 100, -8, -67, -25, 110, 13, 82, -119, -77, -4};
