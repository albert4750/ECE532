wire signed [7:0] convolve1_weight[4][8][3][3];
assign convolve1_weight = '{'{'{'{-1, 116, 3}, '{76, -28, 52}, '{104, -50, 15}}, '{'{20, 99, 58}, '{-105, 79, 13}, '{-11, -43, -80}}, '{'{-79, -59, 41}, '{35, 64, -33}, '{69, -34, -128}}, '{'{-15, 50, -92}, '{34, -80, -35}, '{3, -30, -86}}, '{'{77, -16, 103}, '{21, 73, -1}, '{-128, 10, -14}}, '{'{-85, 58, -1}, '{-105, 59, 2}, '{-7, -30, -66}}, '{'{35, 94, -5}, '{67, -46, 46}, '{99, 20, 81}}, '{'{-78, 27, -114}, '{-87, -70, 65}, '{-92, -118, -42}}}, '{'{'{-85, -24, -117}, '{-126, -77, -48}, '{-96, 54, 0}}, '{'{-90, -109, 46}, '{-86, -13, 56}, '{60, 104, -51}}, '{'{-98, -104, -3}, '{-126, -125, -34}, '{98, -21, -115}}, '{'{-16, -88, -56}, '{-109, -33, -56}, '{26, 66, 120}}, '{'{52, -61, 108}, '{-67, -114, -32}, '{-124, 67, 109}}, '{'{11, 124, -42}, '{77, -7, -19}, '{-53, 56, -112}}, '{'{24, 29, 21}, '{-18, -103, 80}, '{60, -7, -10}}, '{'{-11, 61, -45}, '{33, -24, 32}, '{100, 123, 123}}}, '{'{'{-7, -58, 85}, '{-97, -115, -57}, '{56, 24, -49}}, '{'{-87, -110, -88}, '{54, 79, -117}, '{38, -17, -35}}, '{'{121, 1, 95}, '{-10, -84, 88}, '{-3, -104, -61}}, '{'{82, 111, -125}, '{106, 76, 102}, '{-93, 86, 126}}, '{'{61, 69, 87}, '{-85, -96, -117}, '{-24, 84, 10}}, '{'{54, 107, 37}, '{-3, 28, -17}, '{104, -126, -101}}, '{'{83, 89, 23}, '{-75, -77, 46}, '{20, 53, -99}}, '{'{-61, -93, -89}, '{9, -55, -87}, '{23, 3, -82}}}, '{'{'{90, 50, -20}, '{-125, -97, -119}, '{10, -101, 45}}, '{'{71, 39, -67}, '{-43, -31, -84}, '{-94, 34, -40}}, '{'{-95, 5, 104}, '{127, -92, -128}, '{75, -94, 69}}, '{'{-2, 53, 126}, '{-48, 62, 8}, '{61, 1, 81}}, '{'{-16, -93, -8}, '{-37, 40, -12}, '{-92, 48, -103}}, '{'{-61, -25, 124}, '{-93, -14, -98}, '{-99, 113, -95}}, '{'{18, -111, 93}, '{-44, 125, -126}, '{-59, -27, 12}}, '{'{-84, -11, 125}, '{-62, -17, -37}, '{-43, 39, -89}}}};
