localparam bit signed [0:146][7:0] Input0 = '{-26, -53, -11, 56, 43, 24, -47, -107, 94, 18, -65, -39, -99, -91, 49, 40, 113, -22, 95, -25, -117, -72, 117, 63, 14, -96, 65, -7, -11, -63, -92, 122, -103, 76, -56, -78, -116, 24, 19, 67, 10, -121, 52, -36, -114, 72, -82, 99, -93, 81, 23, -67, -11, 53, -116, 45, -121, 122, 47, -18, 39, -34, 19, 106, -19, 50, -63, 43, -46, 78, 123, -39, -27, -8, 56, -56, 50, -94, 90, -117, -20, 11, -24, 36, -2, 49, 76, 81, 95, 74, -80, -54, 11, -35, -94, 74, 76, 113, -89, -16, -118, -126, -7, 111, -53, 46, -77, 116, 41, 122, -37, 3, -112, -65, -64, -115, -90, -124, -125, 19, -47, 16, -2, -57, 24, -117, 22, -68, 91, 2, 8, -56, 89, -90, -76, 97, -40, -65, 21, -124, 31, 115, 75, 37, -121, 22, -4};
