localparam bit signed [0:26][19:0] Output1 = '{-20'd113, 20'd158, -20'd216, 20'd47, -20'd5, 20'd58, 20'd36, -20'd173, -20'd97, 20'd88, -20'd34, 20'd207, -20'd130, 20'd115, 20'd12, -20'd125, -20'd62, -20'd169, -20'd152, -20'd8, 20'd82, -20'd114, 20'd198, -20'd91, -20'd60, 20'd4, -20'd275};
