localparam bit signed [0:10][15:0] Output1 = '{16'd27105, 16'd16511, -16'd27671, -16'd16486, 16'd19279, -16'd18824, 16'd5248, 16'd5228, -16'd19881, 16'd18651, 16'd25941};
