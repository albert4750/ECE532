logic signed [7:0] layer1_weight[24][3][7][7] = '{
    '{
        '{'{44, -81, -11, 64, -61, 123, 67}, '{-25, -119, 83, -107, 114, -92, -41}, '{-58, 88, -40, 12, -70, 65, 102}, '{-89, -41, 46, -40, -47, 37, -103}, '{-51, -56, -119, 20, -13, 80, 115}, '{69, 126, -49, 47, 64, -46, -29}, '{88, 49, 115, -99, 19, 19, 14}},
        '{'{39, -96, 65, -119, 57, -1, -96}, '{-97, 74, 116, 23, 35, 126, 75}, '{-14, 55, -100, -94, 0, 0, 36}, '{-75, 5, -90, 104, 116, -111, -49}, '{4, -23, -86, 58, -97, -8, -127}, '{-63, 103, 41, -71, -93, -26, -9}, '{-117, 46, -46, -37, 0, 14, -29}},
        '{'{-75, 12, -7, 42, -44, 75, -60}, '{-122, 68, -81, -1, 116, 3, 76}, '{-28, 52, 104, -50, 15, 20, 99}, '{58, -105, 79, 13, -11, -43, -80}, '{-79, -59, 41, 35, 64, -33, 69}, '{-34, -128, -15, 50, -92, 34, -80}, '{-35, 3, -30, -86, 77, -16, 103}}
    },
    '{
        '{'{21, 73, -1, -128, 10, -14, -85}, '{58, -1, -105, 59, 2, -7, -30}, '{-66, 35, 94, -5, 67, -46, 46}, '{99, 20, 81, -78, 27, -114, -87}, '{-70, 65, -92, -118, -42, -85, -24}, '{-117, -126, -77, -48, -96, 54, 0}, '{-90, -109, 46, -86, -13, 56, 60}},
        '{'{104, -51, -98, -104, -3, -126, -125}, '{-34, 98, -21, -115, -16, -88, -56}, '{-109, -33, -56, 26, 66, 120, 52}, '{-61, 108, -67, -114, -32, -124, 67}, '{109, 11, 124, -42, 77, -7, -19}, '{-53, 56, -112, 24, 29, 21, -18}, '{-103, 80, 60, -7, -10, -11, 61}},
        '{'{-45, 33, -24, 32, 100, 123, 123}, '{-7, -58, 85, -97, -115, -57, 56}, '{24, -49, -87, -110, -88, 54, 79}, '{-117, 38, -17, -35, 121, 1, 95}, '{-10, -84, 88, -3, -104, -61, 82}, '{111, -125, 106, 76, 102, -93, 86}, '{126, 61, 69, 87, -85, -96, -117}}
    },
    '{
        '{'{-24, 84, 10, 54, 107, 37, -3}, '{28, -17, 104, -126, -101, 83, 89}, '{23, -75, -77, 46, 20, 53, -99}, '{-61, -93, -89, 9, -55, -87, 23}, '{3, -82, 90, 50, -20, -125, -97}, '{-119, 10, -101, 45, 71, 39, -67}, '{-43, -31, -84, -94, 34, -40, -95}},
        '{'{5, 104, 127, -92, -128, 75, -94}, '{69, -2, 53, 126, -48, 62, 8}, '{61, 1, 81, -16, -93, -8, -37}, '{40, -12, -92, 48, -103, -61, -25}, '{124, -93, -14, -98, -99, 113, -95}, '{18, -111, 93, -44, 125, -126, -59}, '{-27, 12, -84, -11, 125, -62, -17}},
        '{'{-37, -43, 39, -89, 75, 22, 30}, '{17, 70, 71, -110, -36, -85, -45}, '{49, -87, -35, 46, 21, 73, -39}, '{114, 96, 91, -55, -100, 107, 81}, '{-23, 58, 0, 86, -65, -112, -22}, '{36, -34, -104, -12, 63, 67, -77}, '{8, 56, -37, -35, -5, 110, -41}}
    },
    '{
        '{'{32, 19, -56, 71, -41, -115, -70}, '{-47, -8, -12, 55, -64, 75, 92}, '{36, -103, -96, 42, -114, 86, -100}, '{-108, 82, -60, -106, 99, -6, -45}, '{7, 72, -67, 13, -123, -128, 8}, '{79, 79, 53, 11, -124, 39, -36}, '{45, -102, -54, -76, 110, 49, 91}},
        '{'{-77, 99, -23, -110, -11, -94, -77}, '{30, 53, -70, 43, -73, 124, 124}, '{-110, 45, -41, 65, -58, 106, -75}, '{-80, -34, -69, -48, 26, -4, 35}, '{-70, 49, -22, 73, -84, -115, -7}, '{-58, -90, 39, 8, -115, 120, 7}, '{80, 120, -106, 120, -49, 89, -120}},
        '{'{99, -122, 81, 71, 84, 89, 66}, '{-68, 16, -72, -14, 109, 23, -104}, '{-124, -28, 108, -79, -41, -98, -74}, '{25, -108, -31, -27, 57, 23, 27}, '{-99, 33, -13, -75, -9, 51, -42}, '{118, -121, -23, 113, 9, 54, 0}, '{-45, -8, 36, 81, 20, -11, 112}}
    },
    '{
        '{'{-125, -2, -86, -63, -108, -92, -60}, '{80, -16, 47, 10, 109, -24, 94}, '{-37, -85, -65, 31, 20, 70, -119}, '{60, -37, -17, 35, -45, -52, -110}, '{-15, -54, 98, 97, 43, 3, 12}, '{100, -70, 1, -15, 0, -89, -104}, '{58, -92, -29, -59, 6, -125, 98}},
        '{'{-7, 40, 60, 33, -100, -60, -102}, '{96, 120, -19, 51, 73, 53, 69}, '{33, 7, -3, -34, -56, 118, -44}, '{7, 67, 85, 91, -20, -61, -26}, '{-44, -57, -45, 95, -128, 5, -37}, '{-21, 30, 73, 83, -121, 21, 101}, '{92, 8, 43, -82, -128, -24, 51}},
        '{'{-90, -39, -54, 115, 98, -5, -41}, '{-32, -45, -102, 78, -96, -13, 70}, '{-31, 44, -69, -71, 50, 45, 105}, '{4, 57, -35, -37, 17, 35, 66}, '{20, 45, 57, 79, -9, 36, -23}, '{62, -124, 113, 114, 77, 30, -19}, '{-41, 98, 35, -55, 90, 55, -102}}
    },
    '{
        '{'{-10, -106, 76, 79, -30, -38, -77}, '{102, -82, 80, -67, 60, -81, 122}, '{-24, 0, 10, 75, 13, -57, -34}, '{-122, 45, 117, 30, -113, 41, 38}, '{-75, 43, -46, 7, 92, -63, 41}, '{-62, -14, -36, -50, 101, 91, 118}, '{-28, 31, 93, 50, 124, 46, -35}},
        '{'{-14, 33, -116, 96, 105, -48, -62}, '{72, 115, -3, 10, -16, 90, 27}, '{56, -8, -63, 64, 69, -40, -94}, '{79, -125, 60, 110, 37, 43, 83}, '{-40, -58, 20, 6, -100, -13, 6}, '{-62, -36, 92, -26, -27, -5, 69}, '{-19, -55, -28, 54, -51, 21, 123}},
        '{'{31, -47, -93, 109, 115, 122, 8}, '{126, -103, -107, 45, 101, 86, 16}, '{25, 110, -9, 37, -1, 1, 5}, '{70, 12, -38, -54, 123, 54, -50}, '{-66, -56, 71, -83, 5, -81, 59}, '{42, 67, 10, 114, -71, 91, -39}, '{3, -3, 78, -46, 69, 58, 4}}
    },
    '{
        '{'{-111, 69, 63, -34, 24, 3, -59}, '{40, 36, -70, 49, 55, 24, 33}, '{18, -31, 78, 113, 7, 53, 107}, '{-82, 112, 116, -1, 33, -47, 29}, '{-116, -10, -82, -10, -96, -94, -13}, '{-41, -4, 25, 46, 114, -21, -76}, '{105, -18, -64, -52, -10, -55, 18}},
        '{'{-124, -121, 3, -80, -52, -91, -12}, '{109, -80, -19, 82, 51, -79, -57}, '{-38, 49, 110, -99, -125, -54, -44}, '{106, -63, -9, -108, 80, -86, 114}, '{-100, 26, -41, 52, -80, 66, -26}, '{-119, -126, -12, -20, 105, -39, -4}, '{-11, -28, -38, -60, -23, -118, -116}},
        '{'{-24, 97, 37, 39, 32, -6, -95}, '{26, -29, 89, -78, -40, 82, -108}, '{94, 28, -56, -110, 25, 24, -89}, '{106, -5, -100, 24, 18, 67, 44}, '{83, -83, -74, -128, 10, 67, 6}, '{91, -29, 57, 70, 19, 34, -78}, '{114, -26, -108, 43, -10, 0, 100}}
    },
    '{
        '{'{-19, -23, 66, 97, 12, -113, -10}, '{-95, 23, 12, 5, -90, -127, -118}, '{-122, -3, -122, -26, 38, -53, -14}, '{-43, -2, -14, 50, -77, -126, -52}, '{29, -119, -13, 72, 5, -12, 53}, '{107, 65, -85, -49, -66, -52, -81}, '{-52, 21, -8, -110, -39, -115, 94}},
        '{'{-36, 108, -23, 85, -122, -28, -80}, '{-88, 26, 30, 5, 15, 63, 101}, '{-91, -69, -15, -33, -32, 112, 80}, '{-96, -66, 10, 12, -35, -64, 29}, '{-38, 103, 22, 19, 5, -92, -45}, '{-1, 100, -123, -36, 76, 26, 113}, '{-45, 12, 102, 7, 52, -48, 29}},
        '{'{-128, 87, 79, -54, 124, 3, -67}, '{-61, 16, -16, 73, -44, -12, 101}, '{127, -72, -66, 56, -80, 17, -11}, '{57, -119, 108, 62, -49, 102, 78}, '{33, 4, 16, 100, -57, -66, -105}, '{-37, -18, -121, 125, -106, -30, 30}, '{118, -48, 27, -81, 111, -14, -117}}
    },
    '{
        '{'{87, -50, 103, -98, -38, -94, -74}, '{-47, 35, -57, -19, -69, -16, 37}, '{-60, 53, -115, -27, -109, -21, -120}, '{-32, 81, 69, -4, -28, 1, 125}, '{29, 5, 80, 102, 120, 40, 22}, '{-98, 127, -109, -124, 20, -22, -54}, '{-5, 67, 86, -68, 101, 122, -35}},
        '{'{41, -88, 60, 81, 51, -88, -69}, '{106, 94, -99, 97, -34, 110, 37}, '{-2, 88, -112, -29, 39, 29, 124}, '{-63, -105, 72, 0, -41, -91, -17}, '{63, 26, 89, -39, 6, 88, 119}, '{79, -27, -87, 17, 80, -16, -85}, '{-18, 69, -10, 19, 111, -106, -19}},
        '{'{11, -117, 33, 7, -9, -102, -80}, '{71, 111, 54, -32, -28, -46, -41}, '{21, 126, -126, -120, -118, -123, -90}, '{38, -28, 65, -11, -69, 36, 5}, '{-123, -90, 35, -40, 49, 79, -44}, '{-14, -119, 119, 4, 49, -104, -34}, '{2, -45, 3, -51, -117, 13, 100}}
    },
    '{
        '{'{-47, 26, 70, 47, -30, -107, 20}, '{42, -6, 57, 17, -27, 89, 116}, '{85, 55, -28, 68, -17, 98, -117}, '{98, -31, 110, 19, -16, -117, 97}, '{-103, -31, -33, -83, -122, -39, -40}, '{109, -90, -77, -112, 23, 90, -125}, '{-38, 46, -6, 29, -126, 5, -7}},
        '{'{71, -113, -50, 35, 52, -25, -10}, '{-121, 51, -26, 121, 51, 29, 55}, '{-15, 11, 67, 77, -6, -73, -40}, '{123, 124, 120, -60, -11, -13, 86}, '{57, -35, -26, 11, 78, -46, 89}, '{108, -125, 37, 7, -99, -50, -117}, '{73, -117, -112, -68, -5, -25, 63}},
        '{'{59, 1, 18, 53, -100, 64, -43}, '{88, -55, 8, 82, 11, 92, -11}, '{51, -47, 55, -113, 3, -22, 88}, '{85, -100, -70, 85, -50, -17, -63}, '{-52, -117, -103, -25, -117, -38, 109}, '{34, 1, 126, 16, -127, -112, -95}, '{-95, 44, 102, -88, -56, 77, -22}}
    },
    '{
        '{'{-45, 114, 32, 23, -60, 31, 22}, '{-64, 101, -97, -49, -45, -113, -77}, '{121, 12, 45, -118, 116, -23, -48}, '{-58, -107, 94, 67, -48, -64, 1}, '{-78, -32, -21, 123, 82, -46, 57}, '{22, -113, 15, -100, -57, -101, 88}, '{-71, -70, 88, 76, -115, 18, -50}},
        '{'{78, -108, -57, 55, -84, 107, 117}, '{-37, -84, -113, 125, -41, 75, -51}, '{126, 29, -33, -18, 82, 4, -100}, '{65, -79, 49, -41, -71, 80, -87}, '{90, 112, 66, 47, -111, -108, 38}, '{-64, 6, 108, 22, -49, -54, 34}, '{40, 38, 118, 21, -94, -11, 32}},
        '{'{42, -1, -84, -29, -87, 121, -25}, '{27, 123, -80, -1, 10, -60, -111}, '{-125, -27, -34, 87, -99, -26, -5}, '{30, 75, 66, 93, -68, 7, 51}, '{116, -55, 87, 64, 112, 17, 40}, '{115, -107, -34, 26, 15, 112, -111}, '{-118, 17, 3, 103, -55, -99, 67}}
    },
    '{
        '{'{71, 80, 98, 4, 61, -38, -28}, '{6, -96, -47, -9, -10, 117, -91}, '{-9, -101, -77, -50, 59, -42, -33}, '{-120, -72, -99, 28, 95, 34, 58}, '{-1, -2, 81, 92, -17, 16, 72}, '{-69, 119, 108, -121, 12, -96, 84}, '{107, -53, 93, -88, -128, 84, -19}},
        '{'{-36, 77, 37, 47, -67, -25, 50}, '{-60, 110, 76, 57, -9, 101, 112}, '{4, -23, -92, -48, 82, 37, 94}, '{-11, 110, -93, 48, 0, -79, 57}, '{-119, -78, 97, 48, 113, -116, 70}, '{-4, 115, 36, -29, -26, -92, -98}, '{-14, 19, 38, 44, -93, -114, -99}},
        '{'{51, -68, 120, -47, -61, -99, 27}, '{3, -95, 117, 51, -10, 27, 100}, '{-72, -107, 39, 106, -54, -99, 113}, '{29, 61, -70, -104, -14, -112, 64}, '{-28, 98, -5, -115, -127, 123, -126}, '{-62, 19, 116, 122, 76, 30, -89}, '{85, -51, 49, -102, -13, 12, 113}}
    },
    '{
        '{'{64, -127, 36, -118, -22, -96, 126}, '{-100, 58, 66, 92, -63, 77, -45}, '{-81, -47, 36, 71, -75, 70, 9}, '{-113, -110, 29, 53, 60, -86, 82}, '{2, -99, 17, -93, -8, -109, 16}, '{-105, 12, -29, -19, 56, 66, -108}, '{3, -47, 44, -90, -86, 74, -91}},
        '{'{-22, -88, -17, -101, 4, 51, 22}, '{37, -93, -98, -121, 88, -40, 111}, '{15, 10, 19, -51, 103, -72, 101}, '{103, 18, 71, -68, -104, 32, -20}, '{-89, -12, -24, -2, -17, -12, 100}, '{106, -112, 52, 90, 104, 80, -82}, '{96, -34, -44, -105, 15, 44, -45}},
        '{'{-9, -73, -30, 27, -83, 98, -47}, '{87, 27, -51, 48, 87, -34, 5}, '{-7, 103, 97, -15, 98, -100, 116}, '{-63, -60, 85, 72, 124, -14, 33}, '{-10, 99, -80, -29, 89, -59, 65}, '{-29, -57, -127, 1, 71, 25, -28}, '{-51, -20, 50, 27, -32, -85, -109}}
    },
    '{
        '{'{-30, -83, -28, -48, -16, 106, -7}, '{43, 67, -120, 83, 46, -64, -12}, '{20, -32, 98, -21, 5, -43, -104}, '{-126, 125, 125, 71, -20, 75, 115}, '{-100, -10, -33, -63, 80, -14, 82}, '{14, -107, -17, -17, 69, -95, -22}, '{2, -101, 104, -9, 19, 15, -57}},
        '{'{108, -99, 35, 97, -80, 49, -48}, '{56, -65, 88, 58, 5, -77, 122}, '{-67, -22, 83, -111, -83, 96, -66}, '{-106, 97, -26, 9, -123, -52, -67}, '{42, 119, 16, -69, -111, 68, -68}, '{25, 14, -19, -67, 53, -47, -99}, '{70, -100, 74, 5, 100, 100, -44}},
        '{'{55, 114, 50, -42, 53, -118, -85}, '{59, 30, -69, 14, 115, 48, -8}, '{-3, -72, 65, -24, 7, 69, 15}, '{-9, 105, -76, -96, -41, 78, 34}, '{-99, -77, 89, 53, -124, 64, -5}, '{26, 84, 5, -6, -40, -111, 68}, '{-72, 32, 113, -47, -56, -55, 100}}
    },
    '{
        '{'{31, -34, -55, -20, 48, 99, 32}, '{-114, -67, -41, 32, -72, 28, 43}, '{-31, 50, -82, -20, -56, 37, -8}, '{-126, -111, 15, 67, -43, 112, 114}, '{-35, -27, -8, 22, 82, -121, -73}, '{49, -102, 120, 4, -19, -39, -102}, '{60, 115, -17, -45, -50, 18, -7}},
        '{'{-32, -37, -92, -26, 20, -1, 108}, '{3, 18, 77, -77, -79, -97, 97}, '{18, -116, -17, 91, 103, -30, -57}, '{-34, -83, 80, -63, -40, -112, -83}, '{-1, 91, 37, 50, 24, 48, 76}, '{-124, 112, 51, 46, -88, 14, 113}, '{10, 27, -50, -26, 13, -124, 86}},
        '{'{-113, -99, 78, 42, 25, 75, 95}, '{91, -106, -18, -85, 84, 55, 125}, '{2, 25, -3, -8, 0, -33, 56}, '{-18, 70, 82, -42, 62, 127, -82}, '{123, -39, 77, 12, -66, -91, 83}, '{31, -9, 28, -69, 120, -45, -88}, '{-24, -7, -39, 111, -99, -100, -76}}
    },
    '{
        '{'{-86, 10, 84, -111, 0, 39, -90}, '{98, 65, -80, 86, -83, -6, 49}, '{-106, 103, 126, -36, -63, -43, -62}, '{-96, 50, -58, -26, 35, 117, 100}, '{23, 115, -6, -46, -26, -39, 110}, '{-49, -15, 27, -43, -127, -119, -13}, '{-47, 11, -64, 119, -61, 121, 61}},
        '{'{-74, -92, 84, -2, -109, 111, 69}, '{84, -3, 62, 68, 41, 80, 16}, '{57, 5, -32, -106, 3, 8, -66}, '{-36, 41, -54, -26, -36, -33, -20}, '{11, 34, -37, -79, -57, 39, -26}, '{-9, -70, -123, -55, -40, 12, 104}, '{97, -69, 78, 109, -113, -124, 22}},
        '{'{52, -62, -57, -19, -56, -123, -89}, '{-49, -49, -87, 89, 22, 89, 89}, '{19, -66, -99, -119, 11, -3, -29}, '{-102, -25, 127, 82, -56, 127, 1}, '{-29, -14, 113, 46, -73, -118, 74}, '{-104, 127, -33, -85, 91, 13, 78}, '{-73, -123, 23, -86, -25, -79, -27}}
    },
    '{
        '{'{-26, -53, -11, 56, 43, 24, -47}, '{-107, 94, 18, -65, -39, -99, -91}, '{49, 40, 113, -22, 95, -25, -117}, '{-72, 117, 63, 14, -96, 65, -7}, '{-11, -63, -92, 122, -103, 76, -56}, '{-78, -116, 24, 19, 67, 10, -121}, '{52, -36, -114, 72, -82, 99, -93}},
        '{'{81, 23, -67, -11, 53, -116, 45}, '{-121, 122, 47, -18, 39, -34, 19}, '{106, -19, 50, -63, 43, -46, 78}, '{123, -39, -27, -8, 56, -56, 50}, '{-94, 90, -117, -20, 11, -24, 36}, '{-2, 49, 76, 81, 95, 74, -80}, '{-54, 11, -35, -94, 74, 76, 113}},
        '{'{-89, -16, -118, -126, -7, 111, -53}, '{46, -77, 116, 41, 122, -37, 3}, '{-112, -65, -64, -115, -90, -124, -125}, '{19, -47, 16, -2, -57, 24, -117}, '{22, -68, 91, 2, 8, -56, 89}, '{-90, -76, 97, -40, -65, 21, -124}, '{31, 115, 75, 37, -121, 22, -4}}
    },
    '{
        '{'{-86, 59, 95, -74, 73, -13, 51}, '{-46, -105, -45, -103, -71, 69, -39}, '{-83, -17, -40, 51, -69, 44, 26}, '{-8, -11, 43, -7, 32, -98, 14}, '{-57, -32, 61, -127, 118, 47, -4}, '{-19, -10, 43, 90, -113, -60, 74}, '{-43, 39, -22, 107, -34, 86, -128}},
        '{'{-47, 58, -116, 91, -85, 54, -3}, '{47, -106, -97, -12, -94, 98, -86}, '{-60, -6, -66, -92, -45, 44, 81}, '{112, -17, 70, -122, 48, 9, -100}, '{-51, 56, 9, 85, -62, -119, -18}, '{120, 36, -100, 116, -64, 74, -4}, '{13, 107, -126, 37, 71, -41, 94}},
        '{'{81, -125, -17, 98, -48, 115, -46}, '{-78, 61, 106, 82, -100, -93, -75}, '{-102, -15, -25, -86, -82, 69, -100}, '{-1, 43, -45, -66, -54, 74, 9}, '{91, 99, -53, -32, 38, -97, 115}, '{22, -2, -37, -71, -107, 97, -67}, '{108, -87, -13, -21, -29, 41, 122}}
    },
    '{
        '{'{23, 125, 104, -76, -105, -6, -56}, '{-87, 109, -68, -81, 15, -92, 65}, '{-34, 101, -86, 126, -128, 83, 6}, '{93, -61, -97, -99, -112, 67, -102}, '{125, -122, 105, 101, -117, -47, -73}, '{-3, -85, -61, -108, 91, 127, -9}, '{92, -114, -114, -48, 99, 63, -11}},
        '{'{102, -85, 27, -26, 87, 20, 123}, '{-105, -94, -96, -63, -106, -107, 57}, '{-60, -83, 104, 39, -104, -42, -111}, '{52, 90, 8, -123, 97, -42, 122}, '{-46, -118, -66, -99, 11, 30, -57}, '{-70, 94, -86, 85, -57, 25, 108}, '{-74, -10, -45, -103, 45, -7, 106}},
        '{'{3, -12, 84, 113, -45, 121, -91}, '{33, 60, -20, 89, -121, 60, 37}, '{-44, 122, -30, -112, 45, 104, 39}, '{-95, -31, -63, 73, -41, -60, -104}, '{-122, -31, -14, 127, -68, 88, -67}, '{116, 59, 119, -7, 74, -99, 111}, '{120, -100, 24, 3, 82, 21, -122}}
    },
    '{
        '{'{-44, -107, -9, -101, 26, 89, 64}, '{-18, 3, -75, -91, -121, -8, -48}, '{75, 11, 108, 2, -74, -123, -111}, '{122, -3, -50, 5, -50, -47, 105}, '{-18, -20, -98, -30, -125, 0, -35}, '{-84, 44, 108, -1, -13, 61, 126}, '{-128, -111, 29, -37, 34, 114, 115}},
        '{'{100, 59, -107, -65, 94, 120, -27}, '{17, -90, 79, 1, 15, 105, 86}, '{109, -111, 108, 53, 22, 77, -14}, '{47, 66, -117, 9, 114, -88, 54}, '{51, -81, -124, 10, 113, 126, 6}, '{-10, 44, -56, 8, 72, 108, 101}, '{-110, -126, 69, 93, 121, 101, -28}},
        '{'{-22, 29, 27, 17, 58, 11, -79}, '{-56, -40, -125, -16, -117, -71, 50}, '{15, 57, 3, -10, 100, 60, 39}, '{126, 85, 29, 53, -61, -72, 75}, '{-9, -49, -83, -38, -49, 97, -117}, '{119, 5, 30, 58, -60, -69, -96}, '{-91, 43, -3, -68, -83, -99, 122}}
    },
    '{
        '{'{27, 103, -101, -99, -2, -56, -53}, '{-31, 78, -90, -117, 74, 118, -39}, '{-96, 50, -88, 70, -98, 22, -5}, '{-53, -93, 84, 68, -65, -124, 49}, '{-12, 29, 63, -67, -37, -17, 83}, '{-24, -38, -102, -55, 50, 95, -34}, '{-111, 71, -72, 115, -93, 73, 92}},
        '{'{-81, -80, -9, 71, -11, -61, -5}, '{71, -66, 72, -91, -123, -31, -73}, '{92, 46, -90, -79, -120, -6, 65}, '{-62, -66, -112, 61, 66, -117, 31}, '{10, -108, -28, -114, -8, -76, 71}, '{29, 5, -114, -14, 110, 79, -77}, '{-96, 23, 121, -37, -122, 73, -8}},
        '{'{-63, -53, -41, 124, 70, -88, 60}, '{-92, 12, 35, -66, 69, -66, 58}, '{-52, -110, 0, -127, 84, 77, -38}, '{-16, -21, 21, -50, -115, 104, -61}, '{-23, 17, -123, -102, 63, 27, 107}, '{109, 41, -115, -83, 48, -72, -70}, '{-111, 86, -33, 89, 92, 77, 7}}
    },
    '{
        '{'{-102, -111, 68, -85, 47, 94, -3}, '{-36, 121, -56, 58, -101, -122, 7}, '{53, -9, 120, -102, -5, 75, -91}, '{-35, 49, -108, 93, -9, 56, 61}, '{55, 92, 23, 57, 9, 0, -26}, '{19, 71, -78, -90, 67, 124, 30}, '{-91, 56, -2, 105, 5, -69, 80}},
        '{'{90, 61, -97, 70, -39, 75, 17}, '{-97, 31, -44, -38, -89, 117, 50}, '{-54, -90, -60, -5, -89, -1, 79}, '{-115, 35, 102, -5, 11, -25, -53}, '{112, -74, 36, -46, 75, 51, 34}, '{58, -48, -100, 9, -27, -120, 17}, '{112, 108, 92, 25, -34, -5, -27}},
        '{'{59, -5, 94, 121, -69, 58, -110}, '{-116, 1, -101, -118, 67, 61, -112}, '{-101, -4, -122, -128, -121, 25, -61}, '{-69, 120, -12, 127, 36, 44, 85}, '{-15, 118, 127, 72, -17, 38, 42}, '{97, 36, -60, -37, -115, 13, 41}, '{-56, 6, -34, 12, -30, 3, 104}}
    },
    '{
        '{'{-112, -123, -88, 55, 29, 53, -106}, '{-27, -105, 123, -6, 36, 107, 59}, '{-94, 70, 6, -40, -52, -111, -33}, '{-80, -91, -128, 74, -15, -20, -124}, '{-33, 60, -1, -118, -99, -31, -23}, '{112, -115, -109, -87, 76, 44, -77}, '{-21, 16, 120, 126, 114, 37, -114}},
        '{'{36, -14, 4, 114, -81, 0, -79}, '{37, 126, 75, -84, -59, -24, 110}, '{-112, -112, -118, -123, 23, 47, -61}, '{38, 112, -110, -34, 80, -97, 42}, '{-81, -107, 97, -73, -54, -20, -97}, '{-45, -62, 19, 31, -14, -109, -89}, '{39, -67, -31, 44, 116, 108, 54}},
        '{'{94, -6, 103, 62, 76, 16, -48}, '{126, 6, 68, -83, 84, 122, 30}, '{-52, -5, 53, 33, -38, 18, 6}, '{-8, 2, 26, 110, -103, -115, 63}, '{91, -66, -71, -91, 45, 21, -21}, '{120, -59, 121, -79, -103, -116, -76}, '{-58, 47, 125, -55, 10, -56, 90}}
    },
    '{
        '{'{16, -33, -34, 126, 101, -90, 48}, '{60, -122, 112, 70, -9, -127, -17}, '{63, 65, -3, -107, -82, -128, 86}, '{36, 26, 20, -44, 103, -94, 113}, '{-18, -67, 30, 27, 100, -55, -56}, '{-76, -44, 23, -66, -80, 103, 59}, '{-85, 42, 13, 120, -17, 121, -119}},
        '{'{27, -38, 101, -94, -58, 41, 109}, '{-91, -122, -70, -43, -125, -53, 106}, '{-117, 29, -50, 83, -102, -21, 127}, '{-48, 35, -76, 17, -48, 10, 121}, '{60, 73, -29, 25, -1, 26, -77}, '{-49, -101, 4, -26, 85, -25, 113}, '{53, -105, 108, 102, -21, -21, -106}},
        '{'{-36, 110, -85, -122, 13, 77, 17}, '{40, -3, 94, 68, -110, 112, 2}, '{-101, 8, 107, 79, -77, 87, 47}, '{-65, 30, -115, -36, 46, 14, 114}, '{46, 45, -31, -124, -12, 10, -12}, '{-65, -110, 100, 72, -9, -70, 73}, '{110, 13, -116, 29, -50, -24, -51}}
    }
};
