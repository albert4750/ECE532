localparam bit signed [0:15][7:0] Output9 = '{-64, -23, 64, -37, 110, -38, 61, -96, 63, 46, -83, 97, -101, -30, 64, -82};
