localparam bit signed [0:10][0:46][15:0] Weight = '{
    '{-16'd30036, 16'd10799, 16'd9845, 16'd19648, 16'd13123, -16'd11525, -16'd2365, -16'd665, 16'd9225, 16'd24275, -16'd12011, 16'd22258, 16'd14116, -16'd17833, -16'd17338, 16'd15832, 16'd6744, 16'd19852, -16'd18118, -16'd15679, -16'd538, -16'd13785, 16'd10327, 16'd18606, -16'd8616, 16'd2897, 16'd26277, -16'd15847, -16'd5299, 16'd6216, -16'd25847, 16'd6036, -16'd30605, -16'd27696, 16'd4851, -16'd24891, -16'd14338, -16'd30897, -16'd25169, -16'd30272, 16'd15186, -16'd8093, 16'd10200, -16'd847, 16'd755, -16'd31971, 16'd17043},
    '{-16'd29549, -16'd17522, -16'd7769, 16'd23840, -16'd16447, 16'd19721, -16'd13639, 16'd21119, 16'd8736, 16'd23071, 16'd17098, -16'd14092, 16'd24727, 16'd27299, -16'd1538, -16'd21045, 16'd11122, -16'd15177, 16'd22556, 16'd25378, 16'd10368, -16'd6016, 16'd26532, -16'd9163, -16'd26747, -16'd12762, -16'd29208, -16'd7436, 16'd28945, -16'd1713, 16'd12676, 16'd18025, 16'd27690, 16'd13754, 16'd14879, -16'd11400, -16'd12031, 16'd30017, -16'd4121, 16'd28585, -16'd6087, -16'd18141, -16'd20634, 16'd27767, 16'd15115, 16'd8622, 16'd23634},
    '{-16'd12197, 16'd30592, 16'd27022, 16'd19043, -16'd22987, -16'd13428, -16'd5511, -16'd16470, -16'd20396, 16'd18635, -16'd28348, 16'd13062, 16'd7108, -16'd15313, 16'd29311, -16'd18444, 16'd5251, 16'd29644, -16'd25756, -16'd23372, 16'd14312, -16'd28850, -16'd23409, 16'd18068, 16'd11491, -16'd9286, -16'd17641, 16'd10959, 16'd2957, 16'd4469, -16'd18603, -16'd24016, 16'd30001, 16'd9797, -16'd18263, -16'd26973, 16'd17856, -16'd9121, 16'd7365, -16'd4514, 16'd8448, 16'd22385, 16'd3762, 16'd29988, 16'd26530, -16'd7376, -16'd16547},
    '{-16'd13949, 16'd1634, 16'd15914, -16'd31795, -16'd11920, -16'd22553, -16'd21611, -16'd7991, 16'd27007, -16'd18944, 16'd30602, -16'd30350, -16'd19925, -16'd19526, 16'd3455, 16'd22551, 16'd22203, 16'd28802, -16'd26247, -16'd10142, 16'd24126, -16'd23645, -16'd1314, 16'd30843, 16'd10179, 16'd23122, -16'd18514, 16'd19171, -16'd9068, 16'd4305, 16'd18994, 16'd5531, -16'd9458, -16'd983, 16'd31802, -16'd17727, 16'd23588, -16'd9462, 16'd4182, 16'd15403, -16'd19608, -16'd6133, 16'd15106, 16'd307, -16'd19376, -16'd18400, -16'd27466},
    '{16'd1152, -16'd9434, 16'd8467, 16'd5294, 16'd13866, 16'd13683, 16'd17592, 16'd2492, -16'd5656, 16'd15949, 16'd14622, -16'd19176, -16'd7555, 16'd770, -16'd16893, -16'd24482, 16'd11490, 16'd5995, 16'd32013, 16'd30576, -16'd14040, -16'd19128, -16'd29677, 16'd12895, -16'd28856, 16'd17818, -16'd26174, -16'd11016, 16'd24756, 16'd26947, -16'd9236, -16'd24771, 16'd20238, 16'd8032, -16'd17148, 16'd8131, -16'd27923, -16'd6005, 16'd21500, 16'd10838, -16'd29235, -16'd29831, -16'd6547, 16'd4939, 16'd31416, 16'd9744, -16'd13160},
    '{-16'd27747, -16'd5995, 16'd1134, 16'd16409, 16'd9680, -16'd15428, -16'd30855, 16'd19318, -16'd19339, 16'd26045, -16'd18861, 16'd2721, -16'd22680, 16'd17312, -16'd17180, 16'd5627, 16'd27387, 16'd22649, 16'd5446, -16'd32299, 16'd10527, -16'd24051, 16'd18247, 16'd1720, 16'd5272, -16'd15793, 16'd6185, 16'd18706, -16'd16856, -16'd4682, -16'd16177, -16'd17653, 16'd20646, -16'd18321, 16'd19805, -16'd4103, 16'd21633, 16'd31455, 16'd10102, -16'd21716, 16'd24792, -16'd17027, 16'd24600, -16'd4029, 16'd11218, -16'd27665, 16'd24323},
    '{16'd2282, -16'd31028, 16'd22502, -16'd20189, -16'd26922, 16'd13310, 16'd15037, -16'd12603, -16'd29993, -16'd13781, -16'd2016, -16'd9205, -16'd18840, -16'd26412, 16'd1162, 16'd14006, -16'd4117, 16'd30117, -16'd16771, 16'd32412, 16'd623, -16'd536, -16'd23806, 16'd30235, -16'd12333, 16'd1241, 16'd10903, 16'd25397, -16'd28365, -16'd15186, -16'd2924, -16'd13387, 16'd5661, -16'd16829, -16'd21981, -16'd15577, 16'd28041, -16'd30647, 16'd12585, 16'd31639, -16'd8317, -16'd28882, 16'd8922, -16'd10318, -16'd17556, -16'd22781, 16'd18207},
    '{16'd15113, 16'd28042, 16'd28187, 16'd12717, -16'd16185, 16'd1447, -16'd27587, 16'd10581, 16'd29537, 16'd27692, -16'd21726, 16'd10146, -16'd27560, -16'd26591, 16'd14981, 16'd30952, -16'd27905, 16'd22564, 16'd18176, 16'd17867, 16'd14626, -16'd24379, -16'd31874, 16'd30645, 16'd21758, 16'd15440, -16'd2626, 16'd136, -16'd5955, 16'd6273, 16'd26833, -16'd6800, 16'd14627, -16'd19080, -16'd29349, -16'd16216, -16'd26764, 16'd2852, 16'd12464, 16'd9753, -16'd11965, 16'd24423, 16'd25084, -16'd17629, 16'd3186, -16'd10466, -16'd11235},
    '{-16'd14607, 16'd19745, 16'd8338, 16'd21777, 16'd20701, -16'd18092, -16'd11779, -16'd30206, -16'd10171, 16'd30053, -16'd7284, 16'd4652, -16'd19595, -16'd5379, 16'd13634, -16'd4497, 16'd22619, -16'd21163, 16'd423, 16'd28199, 16'd32715, -16'd4458, 16'd28062, 16'd28305, 16'd23238, 16'd967, 16'd4370, 16'd9052, -16'd10197, 16'd21587, 16'd433, -16'd19671, -16'd10147, 16'd29870, -16'd14955, 16'd28873, 16'd12121, -16'd13838, -16'd1568, -16'd18469, -16'd16055, -16'd12772, -16'd16405, -16'd7983, 16'd23145, 16'd30650, 16'd3968},
    '{-16'd8234, -16'd449, -16'd31728, -16'd26518, 16'd24740, -16'd7586, -16'd25064, -16'd25996, 16'd5311, 16'd9411, -16'd6861, 16'd12424, -16'd23624, 16'd29531, -16'd5027, 16'd6011, 16'd19182, 16'd29783, 16'd8352, -16'd30573, -16'd28088, 16'd22983, -16'd7081, 16'd19469, -16'd710, 16'd22097, 16'd5240, -16'd22668, 16'd27575, -16'd17600, 16'd10955, 16'd732, 16'd21412, 16'd24857, 16'd13088, -16'd8790, -16'd20722, -16'd11818, -16'd23268, 16'd7444, -16'd46, 16'd19780, 16'd13846, 16'd21731, -16'd9350, 16'd16979, 16'd647},
    '{-16'd20536, -16'd15811, 16'd6797, 16'd5637, 16'd24832, -16'd4984, 16'd11471, 16'd14799, -16'd75, 16'd5259, 16'd9220, 16'd6567, 16'd4444, 16'd19373, 16'd29978, 16'd586, -16'd18636, 16'd21486, -16'd25167, -16'd4901, -16'd21709, -16'd32029, -16'd3223, -16'd11502, -16'd4747, -16'd27358, 16'd15923, 16'd16030, -16'd15947, -16'd28870, -16'd4181, -16'd14537, -16'd23044, 16'd17404, -16'd9454, -16'd31827, -16'd5289, -16'd7743, -16'd21178, 16'd21994, -16'd21451, -16'd23760, -16'd930, -16'd14277, -16'd18096, -16'd6502, -16'd2436}
};
