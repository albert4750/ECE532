logic signed [7:0] convolve13_weight[4][8][3][3] = '{
    '{
        '{'{-37, 92, 103}, '{-21, -25, -29}, '{30, 116, 41}},
        '{'{118, 9, -10}, '{-76, -85, -47}, '{50, 16, -64}},
        '{'{-102, 7, 54}, '{-46, 58, -53}, '{-71, 58, 76}},
        '{'{-115, 72, 104}, '{-110, 17, 42}, '{-84, 98, 75}},
        '{'{-41, -58, 78}, '{-82, -74, 50}, '{-85, -63, 78}},
        '{'{-27, -122, -7}, '{47, 44, -119}, '{-125, 9, -5}},
        '{'{116, 123, -94}, '{94, -127, -90}, '{78, 80, -34}},
        '{'{50, 13, -42}, '{-82, 99, -41}, '{-91, -35, 109}}
    },
    '{
        '{'{106, -38, -46}, '{86, -122, -54}, '{43, -127, 73}},
        '{'{90, 48, -49}, '{17, -109, 126}, '{19, -63, 27}},
        '{'{115, 100, 35}, '{-119, 105, -115}, '{53, -58, 88}},
        '{'{-118, -7, -85}, '{-27, 5, 40}, '{116, -113, -114}},
        '{'{85, -128, -93}, '{-31, 14, -122}, '{-40, 118, -125}},
        '{'{-60, -27, 104}, '{-33, 27, -14}, '{105, -61, -94}},
        '{'{41, -115, -1}, '{-15, 17, -22}, '{40, 109, 74}},
        '{'{-90, -86, -61}, '{-101, 60, 15}, '{114, 34, 100}}
    },
    '{
        '{'{106, -25, 50}, '{-84, -44, -76}, '{25, 75, 44}},
        '{'{-47, 127, 5}, '{-45, 71, 127}, '{-60, -33, -35}},
        '{'{-22, 114, -37}, '{32, 107, 41}, '{82, 29, 13}},
        '{'{114, -20, 9}, '{-74, 8, -103}, '{33, -111, 113}},
        '{'{47, -112, -79}, '{-66, -57, -34}, '{126, 80, -42}},
        '{'{123, 37, -119}, '{46, 12, -40}, '{-3, -11, 22}},
        '{'{56, -50, -83}, '{-95, 62, -124}, '{-59, -3, -52}},
        '{'{41, 12, -128}, '{69, 22, 105}, '{-31, 49, -13}}
    },
    '{
        '{'{-63, 10, 70}, '{-6, -112, 71}, '{27, -90, -21}},
        '{'{-44, 41, 82}, '{-13, 106, 70}, '{38, 34, -15}},
        '{'{74, 127, -25}, '{-88, -88, 27}, '{-34, 123, 36}},
        '{'{-30, -69, -39}, '{27, 56, -1}, '{58, -97, -80}},
        '{'{107, -2, 3}, '{-64, -91, 119}, '{39, -116, -44}},
        '{'{75, -52, -8}, '{-14, 91, 47}, '{-71, 21, -20}},
        '{'{-116, 111, 17}, '{39, 31, -17}, '{29, 55, 65}},
        '{'{-91, -128, -105}, '{13, 8, 84}, '{-75, 82, -48}}
    }
};
