localparam bit signed [0:2][36:0] Bias3 = '{37'd0, 37'd0, 37'd0};
