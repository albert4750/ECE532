localparam bit signed [0:2][0:26][19:0] Input2 = '{
    '{20'd35, 20'd94, -20'd5, 20'd67, -20'd46, 20'd46, 20'd99, 20'd20, 20'd81, -20'd78, 20'd27, -20'd114, -20'd87, -20'd70, 20'd65, -20'd92, -20'd118, -20'd42, -20'd85, -20'd24, -20'd117, -20'd126, -20'd77, -20'd48, -20'd96, 20'd54, 20'd0},
    '{-20'd90, -20'd109, 20'd46, -20'd86, -20'd13, 20'd56, 20'd60, 20'd104, -20'd51, -20'd98, -20'd104, -20'd3, -20'd126, -20'd125, -20'd34, 20'd98, -20'd21, -20'd115, -20'd16, -20'd88, -20'd56, -20'd109, -20'd33, -20'd56, 20'd26, 20'd66, 20'd120},
    '{20'd52, -20'd61, 20'd108, -20'd67, -20'd114, -20'd32, -20'd124, 20'd67, 20'd109, 20'd11, 20'd124, -20'd42, 20'd77, -20'd7, -20'd19, -20'd53, 20'd56, -20'd112, 20'd24, 20'd29, 20'd21, -20'd18, -20'd103, 20'd80, 20'd60, -20'd7, -20'd10}
};
