localparam bit signed [0:2][0:31][0:4][0:4][24:0] Weight3 = '{
    '{'{'{25'd52116, 25'd312698, -25'd990212, 25'd625397, 25'd156349}, '{25'd625397, 25'd1407143, 25'd52116, -25'd104233, 25'd0}, '{25'd625397, 25'd1094444, -25'd625397, -25'd208466, 25'd885979}, '{25'd469048, 25'd729630, -25'd833862, 25'd885979, -25'd677513}, '{25'd573280, -25'd729630, 25'd625397, 25'd1355026, 25'd729630}}, '{'{25'd312698, 25'd1824074, 25'd677513, 25'd260582, 25'd781746}, '{25'd364815, -25'd208466, 25'd729630, -25'd312698, -25'd677513}, '{-25'd312698, -25'd52116, 25'd521164, 25'd885979, -25'd469048}, '{-25'd52116, 25'd208466, -25'd364815, -25'd260582, -25'd156349}, '{-25'd1250794, 25'd1198677, 25'd2084656, 25'd0, -25'd312698}}, '{'{25'd156349, 25'd885979, 25'd1771958, -25'd260582, -25'd1615608}, '{25'd156349, 25'd573280, 25'd1198677, 25'd1876190, -25'd1042328}, '{25'd1094444, 25'd1407143, 25'd2136772, 25'd1250794, 25'd364815}, '{25'd2136772, 25'd2032540, 25'd3126984, 25'd2501587, 25'd52116}, '{25'd1146561, 25'd1511376, 25'd52116, -25'd573280, -25'd1198677}}, '{'{25'd521164, -25'd990212, 25'd52116, -25'd521164, 25'd0}, '{25'd260582, -25'd885979, 25'd260582, -25'd885979, 25'd677513}, '{25'd938095, 25'd156349, 25'd625397, -25'd208466, -25'd416931}, '{25'd521164, 25'd938095, -25'd625397, 25'd833862, -25'd312698}, '{25'd1250794, -25'd573280, -25'd260582, 25'd1511376, 25'd729630}}, '{'{25'd104233, -25'd1511376, 25'd990212, 25'd677513, -25'd1094444}, '{25'd625397, -25'd469048, 25'd521164, 25'd156349, -25'd938095}, '{-25'd416931, -25'd1094444, 25'd364815, 25'd677513, -25'd938095}, '{25'd416931, -25'd208466, -25'd104233, 25'd312698, -25'd364815}, '{25'd208466, 25'd729630, 25'd416931, 25'd1198677, -25'd729630}}, '{'{25'd885979, 25'd156349, 25'd52116, -25'd260582, -25'd2970635}, '{25'd729630, -25'd312698, 25'd573280, -25'd1094444, -25'd3283333}, '{25'd2762169, 25'd1459259, 25'd2241005, 25'd2866402, 25'd1302910}, '{25'd4377777, 25'd4325661, 25'd3596031, 25'd5263756, 25'd3126984}, '{25'd2032540, 25'd0, 25'd2918518, 25'd1928307, -25'd1407143}}, '{'{25'd1667725, 25'd156349, -25'd1198677, -25'd208466, 25'd1355026}, '{25'd729630, -25'd104233, -25'd1667725, -25'd1563492, -25'd156349}, '{25'd1667725, 25'd729630, -25'd1876190, -25'd1250794, 25'd1615608}, '{25'd312698, 25'd312698, -25'd1355026, 25'd833862, 25'd990212}, '{25'd1719841, -25'd469048, 25'd781746, 25'd52116, -25'd364815}}, '{'{25'd1719841, 25'd781746, 25'd1771958, 25'd1719841, -25'd1771958}, '{25'd781746, 25'd2345238, 25'd3126984, 25'd729630, 25'd208466}, '{25'd2188889, 25'd2188889, 25'd3908730, 25'd1876190, 25'd1094444}, '{25'd469048, 25'd1459259, 25'd3231217, 25'd1511376, -25'd1719841}, '{25'd52116, 25'd104233, 25'd2084656, 25'd312698, -25'd1094444}}, '{'{-25'd364815, -25'd990212, 25'd781746, 25'd0, 25'd156349}, '{25'd312698, 25'd260582, 25'd573280, 25'd677513, 25'd0}, '{-25'd781746, -25'd52116, -25'd1042328, -25'd729630, -25'd1042328}, '{25'd625397, 25'd833862, 25'd938095, 25'd416931, 25'd1250794}, '{-25'd469048, 25'd1042328, 25'd1146561, 25'd990212, 25'd1042328}}, '{'{25'd1459259, 25'd1407143, 25'd938095, -25'd104233, 25'd469048}, '{-25'd729630, 25'd416931, 25'd364815, 25'd885979, -25'd833862}, '{25'd573280, 25'd312698, 25'd521164, -25'd885979, 25'd573280}, '{-25'd729630, -25'd104233, 25'd833862, 25'd416931, 25'd885979}, '{25'd1407143, -25'd729630, -25'd1042328, 25'd625397, 25'd364815}}, '{'{-25'd312698, 25'd1355026, 25'd1146561, -25'd833862, 25'd677513}, '{25'd833862, 25'd885979, -25'd573280, 25'd469048, 25'd625397}, '{25'd104233, -25'd781746, 25'd1302910, 25'd1042328, -25'd1042328}, '{25'd885979, 25'd416931, 25'd729630, -25'd1042328, -25'd885979}, '{25'd833862, 25'd1407143, 25'd1094444, -25'd677513, -25'd990212}}, '{'{25'd1980423, -25'd990212, -25'd312698, 25'd312698, 25'd938095}, '{-25'd469048, -25'd1459259, -25'd2032540, -25'd1302910, 25'd1459259}, '{25'd156349, -25'd208466, -25'd1042328, 25'd0, 25'd1928307}, '{25'd573280, -25'd885979, 25'd208466, 25'd260582, 25'd625397}, '{25'd469048, -25'd156349, -25'd260582, 25'd2032540, 25'd1511376}}, '{'{-25'd2188889, 25'd990212, 25'd1146561, -25'd416931, -25'd1407143}, '{25'd208466, 25'd1771958, 25'd1980423, -25'd416931, -25'd3283333}, '{-25'd729630, 25'd729630, 25'd1928307, -25'd260582, -25'd2449471}, '{-25'd729630, 25'd1146561, 25'd2918518, -25'd1459259, -25'd1980423}, '{-25'd2032540, 25'd1511376, 25'd1198677, -25'd1928307, -25'd3439682}}, '{'{-25'd781746, -25'd990212, -25'd1563492, 25'd312698, -25'd573280}, '{25'd156349, -25'd625397, -25'd156349, -25'd1355026, -25'd1459259}, '{-25'd52116, -25'd573280, -25'd1198677, -25'd1302910, 25'd625397}, '{-25'd1302910, 25'd208466, -25'd52116, 25'd573280, 25'd104233}, '{25'd416931, -25'd1302910, -25'd104233, -25'd833862, 25'd1042328}}, '{'{25'd260582, -25'd521164, 25'd364815, 25'd156349, 25'd312698}, '{25'd156349, 25'd1042328, -25'd833862, -25'd677513, -25'd469048}, '{25'd1094444, 25'd521164, 25'd1302910, 25'd729630, 25'd938095}, '{-25'd208466, -25'd260582, -25'd469048, 25'd0, -25'd677513}, '{-25'd260582, 25'd573280, 25'd573280, 25'd625397, 25'd1042328}}, '{'{25'd833862, 25'd1198677, 25'd1042328, 25'd156349, 25'd156349}, '{25'd833862, -25'd104233, -25'd469048, -25'd104233, 25'd990212}, '{-25'd208466, 25'd52116, -25'd208466, 25'd1511376, 25'd1250794}, '{-25'd208466, 25'd1250794, -25'd469048, 25'd521164, 25'd625397}, '{25'd625397, -25'd364815, 25'd990212, -25'd260582, 25'd781746}}, '{'{25'd1667725, -25'd156349, -25'd2032540, 25'd3804497, 25'd2345238}, '{25'd990212, -25'd2084656, -25'd3804497, 25'd416931, 25'd677513}, '{25'd2918518, 25'd260582, -25'd4377777, 25'd833862, 25'd1198677}, '{25'd2970635, 25'd208466, -25'd4012963, 25'd1928307, 25'd1876190}, '{25'd938095, 25'd1250794, -25'd1302910, 25'd1824074, -25'd260582}}, '{'{-25'd521164, 25'd1094444, 25'd469048, -25'd208466, -25'd677513}, '{-25'd677513, 25'd156349, 25'd1094444, -25'd1094444, -25'd156349}, '{-25'd885979, -25'd885979, 25'd885979, -25'd416931, -25'd990212}, '{25'd1146561, -25'd677513, -25'd625397, -25'd1146561, 25'd0}, '{-25'd52116, -25'd469048, 25'd104233, -25'd156349, -25'd364815}}, '{'{25'd2084656, -25'd364815, -25'd729630, 25'd0, 25'd677513}, '{25'd104233, 25'd104233, -25'd1876190, -25'd1980423, 25'd1407143}, '{25'd1667725, 25'd885979, -25'd1198677, -25'd885979, 25'd156349}, '{25'd1198677, -25'd1094444, -25'd990212, 25'd1146561, 25'd104233}, '{-25'd52116, -25'd104233, 25'd1459259, 25'd1250794, 25'd469048}}, '{'{25'd833862, 25'd469048, -25'd625397, 25'd364815, 25'd364815}, '{25'd0, 25'd938095, 25'd0, -25'd364815, 25'd521164}, '{-25'd781746, 25'd1302910, 25'd781746, 25'd156349, 25'd677513}, '{25'd729630, -25'd833862, 25'd52116, 25'd0, 25'd781746}, '{-25'd208466, 25'd260582, 25'd1250794, -25'd1042328, -25'd885979}}, '{'{25'd1146561, 25'd625397, 25'd625397, -25'd573280, -25'd156349}, '{-25'd364815, 25'd781746, -25'd364815, 25'd0, 25'd885979}, '{-25'd990212, 25'd729630, 25'd625397, 25'd260582, -25'd833862}, '{25'd625397, 25'd156349, -25'd312698, -25'd260582, 25'd1042328}, '{25'd990212, -25'd156349, -25'd625397, -25'd312698, -25'd990212}}, '{'{25'd1511376, -25'd625397, 25'd52116, -25'd312698, -25'd156349}, '{25'd1719841, 25'd1511376, 25'd364815, -25'd156349, -25'd208466}, '{-25'd729630, -25'd260582, -25'd52116, -25'd729630, 25'd833862}, '{-25'd312698, 25'd156349, -25'd260582, 25'd104233, 25'd1667725}, '{-25'd573280, -25'd104233, 25'd625397, 25'd104233, 25'd1198677}}, '{'{-25'd2084656, -25'd2241005, 25'd3856613, 25'd4482010, -25'd1876190}, '{25'd416931, 25'd1407143, 25'd4951058, 25'd5472222, -25'd521164}, '{-25'd1719841, -25'd521164, 25'd3543915, 25'd4429894, -25'd2970635}, '{-25'd2397354, -25'd3596031, 25'd1094444, 25'd1302910, -25'd4742592}, '{-25'd2866402, -25'd3126984, -25'd469048, 25'd781746, -25'd4012963}}, '{'{-25'd1771958, -25'd2553704, 25'd521164, -25'd729630, -25'd2032540}, '{-25'd416931, -25'd781746, 25'd677513, -25'd677513, -25'd1615608}, '{25'd2032540, 25'd2084656, 25'd1876190, 25'd1459259, 25'd625397}, '{25'd2084656, 25'd1928307, 25'd3231217, 25'd2397354, 25'd0}, '{25'd1719841, 25'd364815, 25'd3074867, 25'd2136772, -25'd521164}}, '{'{-25'd781746, 25'd208466, -25'd104233, 25'd0, -25'd729630}, '{25'd1459259, 25'd833862, 25'd364815, 25'd1302910, -25'd990212}, '{-25'd938095, -25'd885979, 25'd938095, 25'd104233, -25'd729630}, '{25'd208466, 25'd364815, -25'd416931, 25'd312698, -25'd416931}, '{25'd1511376, 25'd52116, 25'd677513, 25'd677513, -25'd364815}}, '{'{-25'd2032540, -25'd2084656, -25'd260582, -25'd781746, -25'd1094444}, '{25'd104233, -25'd1511376, -25'd52116, -25'd677513, -25'd2501587}, '{-25'd1094444, 25'd416931, 25'd1407143, 25'd573280, -25'd2241005}, '{-25'd2241005, -25'd1042328, 25'd0, -25'd1407143, -25'd1876190}, '{-25'd312698, 25'd0, -25'd1459259, -25'd1042328, -25'd1511376}}, '{'{25'd416931, -25'd208466, 25'd260582, 25'd104233, 25'd781746}, '{25'd729630, 25'd833862, -25'd52116, -25'd573280, 25'd573280}, '{25'd1094444, -25'd260582, -25'd1042328, 25'd1302910, -25'd416931}, '{25'd312698, -25'd990212, 25'd1042328, 25'd104233, -25'd104233}, '{25'd1250794, 25'd416931, -25'd729630, -25'd677513, -25'd729630}}, '{'{25'd1459259, 25'd1250794, -25'd469048, 25'd1146561, 25'd625397}, '{25'd885979, 25'd416931, -25'd260582, 25'd1250794, 25'd52116}, '{-25'd156349, 25'd781746, -25'd781746, -25'd521164, 25'd521164}, '{-25'd208466, -25'd677513, -25'd938095, 25'd364815, -25'd104233}, '{25'd312698, 25'd573280, -25'd260582, -25'd416931, -25'd1042328}}, '{'{-25'd1094444, 25'd416931, 25'd52116, 25'd208466, 25'd364815}, '{-25'd312698, 25'd156349, -25'd1042328, 25'd1198677, -25'd208466}, '{25'd1198677, -25'd625397, -25'd677513, -25'd416931, -25'd781746}, '{25'd885979, 25'd938095, 25'd833862, -25'd885979, -25'd625397}, '{25'd1042328, -25'd469048, -25'd938095, -25'd1042328, -25'd1094444}}, '{'{25'd677513, -25'd469048, 25'd469048, 25'd833862, 25'd677513}, '{25'd573280, -25'd990212, 25'd1042328, 25'd1719841, 25'd1302910}, '{-25'd1094444, 25'd990212, 25'd1094444, 25'd573280, -25'd833862}, '{-25'd52116, -25'd312698, 25'd0, -25'd469048, -25'd521164}, '{25'd1302910, -25'd833862, 25'd364815, 25'd364815, 25'd1042328}}, '{'{-25'd1302910, 25'd104233, 25'd990212, 25'd781746, -25'd3856613}, '{-25'd156349, 25'd364815, 25'd2032540, 25'd2397354, -25'd1302910}, '{25'd625397, -25'd677513, 25'd677513, 25'd2605820, 25'd2397354}, '{-25'd1667725, -25'd2762169, -25'd885979, 25'd1094444, -25'd833862}, '{-25'd2032540, -25'd625397, -25'd1042328, 25'd1771958, 25'd1719841}}, '{'{-25'd2136772, -25'd1615608, -25'd729630, -25'd156349, 25'd1042328}, '{-25'd1250794, -25'd1146561, -25'd1824074, 25'd1042328, -25'd1928307}, '{25'd521164, 25'd2345238, 25'd2553704, 25'd2657936, 25'd1355026}, '{25'd2188889, 25'd1719841, 25'd2657936, 25'd2918518, -25'd2345238}, '{25'd156349, 25'd2136772, 25'd2241005, -25'd2553704, -25'd6670899}}},
    '{'{'{25'd307187, -25'd614375, 25'd716771, -25'd409583, -25'd614375}, '{-25'd1126354, -25'd1228750, -25'd1126354, -25'd614375, 25'd1126354}, '{25'd409583, 25'd614375, 25'd614375, 25'd307187, -25'd614375}, '{25'd1126354, 25'd511979, 25'd1228750, -25'd102396, -25'd716771}, '{25'd307187, -25'd1331146, 25'd102396, -25'd819166, 25'd1126354}}, '{'{-25'd204792, 25'd0, 25'd102396, 25'd1126354, 25'd819166}, '{-25'd204792, 25'd1740729, 25'd1535937, 25'd1843125, 25'd716771}, '{25'd921562, -25'd614375, -25'd511979, 25'd716771, 25'd1023958}, '{25'd102396, -25'd614375, 25'd409583, 25'd819166, -25'd614375}, '{-25'd204792, -25'd511979, -25'd307187, 25'd819166, 25'd1126354}}, '{'{25'd1433541, 25'd0, 25'd1433541, 25'd1433541, -25'd1331146}, '{25'd1023958, 25'd1843125, 25'd3481457, 25'd2150312, -25'd614375}, '{25'd1638333, 25'd2150312, 25'd2150312, 25'd2969478, 25'd2355104}, '{25'd2559895, 25'd3481457, 25'd2047916, 25'd1331146, 25'd1023958}, '{25'd2252708, 25'd2764687, 25'd1023958, 25'd819166, 25'd409583}}, '{'{25'd716771, 25'd1228750, 25'd819166, -25'd204792, 25'd921562}, '{25'd1023958, -25'd204792, 25'd409583, 25'd921562, 25'd204792}, '{-25'd102396, 25'd102396, -25'd307187, -25'd1023958, 25'd511979}, '{25'd1228750, -25'd1228750, 25'd921562, 25'd614375, 25'd614375}, '{25'd204792, 25'd819166, -25'd1126354, -25'd204792, -25'd1126354}}, '{'{-25'd204792, 25'd1126354, 25'd204792, -25'd1331146, 25'd1331146}, '{25'd409583, -25'd1023958, -25'd409583, -25'd1023958, -25'd409583}, '{25'd819166, -25'd614375, 25'd409583, 25'd1023958, -25'd409583}, '{-25'd204792, -25'd409583, -25'd1126354, 25'd409583, -25'd409583}, '{-25'd307187, 25'd1126354, 25'd716771, -25'd511979, 25'd1023958}}, '{'{25'd1945520, 25'd1126354, -25'd1126354, -25'd409583, -25'd1638333}, '{25'd716771, -25'd1843125, -25'd1945520, -25'd2252708, -25'd2252708}, '{25'd1638333, 25'd102396, 25'd1228750, 25'd1843125, -25'd409583}, '{25'd921562, -25'd614375, 25'd1331146, 25'd3686249, 25'd204792}, '{25'd1228750, -25'd409583, 25'd307187, 25'd1843125, -25'd2047916}}, '{'{-25'd204792, -25'd716771, 25'd0, -25'd307187, 25'd1945520}, '{25'd1535937, 25'd614375, -25'd716771, -25'd1023958, 25'd716771}, '{25'd819166, 25'd102396, -25'd307187, -25'd307187, 25'd1740729}, '{25'd1023958, -25'd614375, 25'd716771, 25'd307187, 25'd614375}, '{25'd307187, 25'd1843125, -25'd204792, 25'd1228750, 25'd511979}}, '{'{25'd1023958, 25'd0, 25'd2867083, 25'd1638333, -25'd2662291}, '{25'd1535937, 25'd1740729, 25'd4300624, 25'd2764687, -25'd1535937}, '{25'd1945520, 25'd3276666, 25'd4914999, 25'd1535937, -25'd1535937}, '{25'd1535937, 25'd716771, 25'd3174270, 25'd0, -25'd2457499}, '{-25'd1740729, -25'd1023958, 25'd1126354, -25'd204792, -25'd3891041}}, '{'{-25'd921562, -25'd819166, 25'd0, -25'd921562, 25'd204792}, '{-25'd102396, -25'd409583, 25'd307187, 25'd307187, 25'd0}, '{25'd1023958, 25'd614375, 25'd1228750, -25'd1023958, 25'd921562}, '{25'd409583, 25'd1023958, 25'd921562, -25'd716771, 25'd307187}, '{-25'd614375, -25'd819166, 25'd102396, -25'd1023958, -25'd614375}}, '{'{-25'd716771, 25'd0, -25'd511979, 25'd1228750, -25'd1126354}, '{25'd409583, -25'd1023958, -25'd1126354, -25'd307187, -25'd204792}, '{25'd1228750, 25'd921562, 25'd819166, -25'd614375, 25'd204792}, '{25'd819166, -25'd614375, -25'd1126354, 25'd1228750, 25'd921562}, '{-25'd511979, 25'd1331146, 25'd307187, -25'd511979, -25'd511979}}, '{'{-25'd409583, -25'd614375, -25'd204792, -25'd307187, -25'd102396}, '{25'd1023958, -25'd204792, 25'd409583, -25'd409583, 25'd1331146}, '{25'd511979, 25'd409583, 25'd819166, -25'd1023958, -25'd1126354}, '{-25'd409583, -25'd1228750, 25'd1023958, 25'd1023958, -25'd716771}, '{25'd511979, 25'd102396, 25'd307187, 25'd0, 25'd511979}}, '{'{25'd2047916, -25'd614375, -25'd2355104, -25'd1126354, 25'd2150312}, '{25'd1433541, -25'd2150312, -25'd2047916, -25'd716771, 25'd1023958}, '{25'd819166, -25'd2047916, -25'd409583, -25'd409583, 25'd2559895}, '{25'd1945520, -25'd1331146, 25'd819166, 25'd2150312, 25'd1945520}, '{-25'd102396, 25'd614375, -25'd716771, 25'd1433541, 25'd1843125}}, '{'{-25'd3071874, -25'd1126354, 25'd102396, -25'd1433541, -25'd1331146}, '{-25'd1638333, 25'd1228750, 25'd1331146, -25'd1126354, -25'd1023958}, '{-25'd1740729, 25'd204792, 25'd716771, -25'd1740729, -25'd2457499}, '{-25'd2355104, -25'd102396, 25'd1535937, -25'd1023958, -25'd2559895}, '{-25'd1945520, -25'd102396, 25'd1331146, -25'd1638333, -25'd2662291}}, '{'{-25'd1126354, 25'd102396, -25'd1126354, -25'd409583, -25'd921562}, '{-25'd1023958, -25'd1228750, 25'd1023958, -25'd921562, 25'd614375}, '{-25'd1331146, -25'd1023958, 25'd511979, 25'd921562, 25'd1126354}, '{25'd614375, 25'd307187, -25'd614375, 25'd614375, 25'd102396}, '{-25'd1023958, -25'd1023958, -25'd1126354, -25'd921562, -25'd716771}}, '{'{-25'd204792, 25'd307187, -25'd102396, -25'd307187, 25'd1228750}, '{-25'd307187, 25'd409583, -25'd614375, -25'd1228750, 25'd819166}, '{25'd614375, 25'd1126354, -25'd307187, 25'd204792, 25'd1023958}, '{25'd1228750, 25'd1331146, -25'd409583, 25'd716771, 25'd1023958}, '{25'd716771, 25'd1228750, 25'd307187, 25'd716771, 25'd716771}}, '{'{25'd409583, 25'd921562, -25'd204792, -25'd409583, 25'd307187}, '{25'd716771, 25'd921562, 25'd921562, -25'd204792, 25'd716771}, '{-25'd307187, 25'd614375, 25'd0, 25'd819166, 25'd921562}, '{-25'd102396, 25'd102396, -25'd409583, -25'd204792, 25'd409583}, '{25'd0, -25'd921562, -25'd1433541, -25'd1331146, 25'd307187}}, '{'{25'd1638333, 25'd0, -25'd3993437, 25'd2355104, 25'd2150312}, '{-25'd2355104, -25'd2764687, -25'd7065311, -25'd3993437, -25'd1638333}, '{-25'd307187, -25'd511979, -25'd5734165, 25'd614375, 25'd1126354}, '{25'd614375, 25'd511979, -25'd4710207, 25'd2457499, 25'd4300624}, '{25'd511979, 25'd2355104, -25'd4607811, 25'd2867083, 25'd3891041}}, '{'{25'd1843125, 25'd0, 25'd1843125, 25'd102396, -25'd1023958}, '{25'd1843125, -25'd409583, 25'd0, 25'd409583, 25'd1228750}, '{-25'd409583, 25'd307187, 25'd0, -25'd307187, -25'd819166}, '{-25'd614375, 25'd1433541, 25'd409583, 25'd921562, 25'd614375}, '{-25'd1023958, -25'd102396, -25'd819166, 25'd921562, 25'd307187}}, '{'{25'd1638333, 25'd716771, -25'd1023958, 25'd102396, 25'd1740729}, '{25'd1740729, -25'd1023958, -25'd1023958, -25'd614375, 25'd614375}, '{25'd0, -25'd204792, -25'd204792, -25'd1023958, 25'd819166}, '{25'd1023958, 25'd102396, 25'd921562, 25'd409583, -25'd819166}, '{25'd0, -25'd409583, 25'd921562, 25'd102396, 25'd511979}}, '{'{25'd0, 25'd1126354, -25'd409583, 25'd1023958, 25'd1331146}, '{25'd1126354, -25'd511979, -25'd1023958, -25'd511979, 25'd307187}, '{25'd819166, -25'd614375, 25'd204792, -25'd511979, 25'd102396}, '{25'd819166, 25'd921562, 25'd511979, -25'd307187, 25'd102396}, '{25'd409583, 25'd102396, 25'd614375, 25'd819166, 25'd819166}}, '{'{25'd1126354, 25'd819166, 25'd921562, 25'd511979, -25'd819166}, '{25'd614375, -25'd1023958, -25'd614375, 25'd614375, 25'd204792}, '{25'd921562, 25'd0, 25'd1331146, -25'd204792, -25'd1126354}, '{25'd614375, -25'd819166, 25'd1023958, 25'd819166, 25'd1023958}, '{25'd716771, 25'd511979, 25'd716771, -25'd1126354, 25'd0}}, '{'{25'd614375, 25'd204792, 25'd102396, -25'd511979, -25'd819166}, '{25'd1228750, 25'd1331146, 25'd819166, -25'd716771, 25'd1228750}, '{25'd1331146, 25'd102396, -25'd614375, -25'd307187, 25'd409583}, '{25'd102396, -25'd614375, -25'd307187, 25'd409583, 25'd511979}, '{25'd1331146, 25'd921562, -25'd819166, 25'd307187, 25'd1331146}}, '{'{-25'd1638333, -25'd1638333, 25'd2867083, 25'd3174270, 25'd511979}, '{-25'd1535937, 25'd819166, 25'd3276666, 25'd3481457, -25'd204792}, '{-25'd3174270, -25'd1126354, 25'd2150312, 25'd1740729, -25'd1843125}, '{-25'd3379062, -25'd1331146, -25'd1331146, 25'd0, -25'd2150312}, '{-25'd2559895, -25'd2047916, 25'd1740729, -25'd102396, -25'd3276666}}, '{'{-25'd1843125, -25'd1740729, 25'd307187, -25'd511979, -25'd2969478}, '{-25'd307187, -25'd1535937, -25'd614375, -25'd1228750, -25'd307187}, '{25'd1331146, 25'd921562, 25'd716771, 25'd2457499, -25'd614375}, '{25'd716771, 25'd511979, 25'd1843125, 25'd307187, -25'd614375}, '{-25'd1638333, 25'd1228750, 25'd614375, -25'd102396, -25'd1228750}}, '{'{-25'd819166, 25'd1023958, -25'd614375, 25'd307187, -25'd511979}, '{25'd716771, -25'd204792, 25'd614375, 25'd0, 25'd921562}, '{25'd819166, 25'd614375, 25'd1228750, 25'd1023958, -25'd102396}, '{25'd1228750, 25'd716771, 25'd1228750, -25'd102396, 25'd511979}, '{-25'd614375, -25'd409583, 25'd204792, 25'd1023958, -25'd819166}}, '{'{25'd409583, 25'd102396, 25'd2047916, 25'd511979, 25'd0}, '{25'd511979, 25'd2764687, 25'd3379062, 25'd1740729, 25'd0}, '{25'd614375, 25'd1638333, 25'd2662291, 25'd2047916, 25'd819166}, '{25'd921562, 25'd1126354, 25'd3481457, 25'd1638333, 25'd716771}, '{25'd2252708, 25'd2867083, 25'd3174270, 25'd1945520, 25'd1638333}}, '{'{25'd1023958, -25'd614375, 25'd409583, -25'd204792, 25'd1023958}, '{-25'd819166, -25'd511979, 25'd716771, -25'd921562, -25'd921562}, '{25'd204792, -25'd1126354, 25'd1023958, -25'd511979, 25'd819166}, '{-25'd307187, 25'd614375, 25'd204792, -25'd1126354, -25'd921562}, '{25'd819166, 25'd307187, -25'd819166, 25'd511979, 25'd819166}}, '{'{-25'd716771, 25'd409583, -25'd819166, 25'd819166, 25'd716771}, '{-25'd921562, 25'd1126354, -25'd716771, 25'd0, -25'd921562}, '{25'd614375, 25'd614375, -25'd819166, -25'd819166, -25'd716771}, '{25'd716771, 25'd307187, 25'd0, 25'd1228750, 25'd409583}, '{25'd1126354, 25'd1023958, 25'd511979, -25'd819166, 25'd1126354}}, '{'{25'd716771, 25'd716771, 25'd0, 25'd307187, 25'd614375}, '{-25'd921562, -25'd409583, -25'd511979, 25'd102396, -25'd511979}, '{-25'd409583, 25'd614375, 25'd409583, 25'd1023958, 25'd1228750}, '{-25'd1126354, -25'd1023958, -25'd921562, -25'd1023958, -25'd614375}, '{25'd511979, -25'd409583, -25'd819166, -25'd307187, -25'd716771}}, '{'{25'd511979, -25'd716771, 25'd0, 25'd1638333, 25'd819166}, '{25'd921562, -25'd614375, 25'd716771, 25'd1638333, 25'd1228750}, '{25'd1228750, 25'd1126354, 25'd1331146, 25'd511979, 25'd614375}, '{-25'd204792, 25'd511979, -25'd819166, 25'd0, -25'd716771}, '{25'd102396, 25'd409583, 25'd0, -25'd819166, 25'd102396}}, '{'{-25'd1740729, -25'd1740729, 25'd1331146, 25'd921562, -25'd7986873}, '{25'd1433541, 25'd2252708, 25'd2252708, 25'd2252708, 25'd2252708}, '{25'd511979, 25'd409583, 25'd1740729, 25'd3481457, 25'd3276666}, '{-25'd1023958, -25'd1535937, 25'd409583, 25'd1023958, 25'd819166}, '{-25'd1228750, 25'd204792, -25'd511979, 25'd1638333, 25'd0}}, '{'{25'd102396, -25'd1740729, -25'd2559895, 25'd921562, -25'd1228750}, '{25'd204792, -25'd921562, -25'd1126354, 25'd1843125, -25'd614375}, '{25'd3071874, 25'd1945520, 25'd3788645, 25'd4812603, 25'd614375}, '{25'd2150312, 25'd4505416, 25'd4198228, 25'd5017395, -25'd3071874}, '{-25'd2867083, 25'd1228750, 25'd1228750, -25'd4914999, -25'd13106663}}},
    '{'{'{-25'd901062, 25'd732113, 25'd506847, -25'd844746, -25'd619480}, '{-25'd168949, 25'd1182644, 25'd225266, 25'd0, 25'd675797}, '{25'd394215, -25'd957378, -25'd619480, -25'd112633, 25'd957378}, '{-25'd957378, 25'd168949, -25'd957378, 25'd56316, -25'd732113}, '{25'd957378, -25'd1182644, 25'd337898, 25'd225266, -25'd675797}}, '{'{25'd281582, 25'd394215, 25'd901062, 25'd957378, 25'd1858441}, '{-25'd56316, 25'd901062, 25'd563164, 25'd450531, -25'd56316}, '{-25'd1126328, -25'd563164, 25'd1633175, 25'd1351593, -25'd168949}, '{25'd394215, 25'd844746, -25'd225266, 25'd1407909, 25'd1013695}, '{-25'd56316, -25'd450531, 25'd225266, 25'd1182644, 25'd563164}}, '{'{25'd0, 25'd281582, 25'd1013695, -25'd619480, -25'd1013695}, '{25'd1126328, 25'd1295277, 25'd1013695, 25'd394215, -25'd732113}, '{25'd1576859, 25'd619480, 25'd675797, 25'd2646870, -25'd281582}, '{25'd732113, 25'd2759503, 25'd844746, 25'd788429, 25'd1295277}, '{25'd281582, 25'd1351593, 25'd1633175, 25'd1576859, -25'd1295277}}, '{'{-25'd788429, 25'd675797, -25'd168949, 25'd901062, 25'd788429}, '{25'd0, 25'd901062, -25'd563164, 25'd957378, 25'd732113}, '{-25'd901062, -25'd225266, -25'd675797, -25'd675797, 25'd1238960}, '{25'd732113, -25'd56316, 25'd225266, -25'd844746, 25'd901062}, '{-25'd1013695, 25'd56316, 25'd1070011, -25'd563164, 25'd0}}, '{'{-25'd732113, 25'd957378, -25'd225266, 25'd337898, -25'd1182644}, '{25'd1295277, 25'd1295277, 25'd0, -25'd788429, -25'd619480}, '{-25'd506847, -25'd788429, 25'd1576859, -25'd619480, 25'd56316}, '{-25'd506847, -25'd506847, 25'd1295277, -25'd563164, 25'd450531}, '{25'd281582, 25'd675797, 25'd675797, -25'd1013695, -25'd563164}}, '{'{25'd2140022, 25'd168949, -25'd2477921, -25'd1914757, -25'd732113}, '{25'd56316, -25'd1295277, -25'd1464226, -25'd1520542, -25'd1914757}, '{25'd2083706, -25'd1126328, -25'd957378, 25'd2984768, 25'd112633}, '{25'd1070011, -25'd675797, -25'd2083706, -25'd168949, -25'd2759503}, '{25'd1295277, -25'd1182644, -25'd732113, 25'd1070011, -25'd337898}}, '{'{25'd2027390, 25'd732113, -25'd1295277, -25'd1070011, 25'd1576859}, '{25'd901062, 25'd450531, -25'd1745808, -25'd844746, 25'd1689491}, '{25'd225266, 25'd1126328, -25'd563164, -25'd957378, 25'd56316}, '{25'd1745808, 25'd675797, -25'd1407909, 25'd901062, 25'd337898}, '{25'd1802124, 25'd563164, 25'd1295277, 25'd1182644, -25'd1013695}}, '{'{-25'd56316, -25'd1013695, 25'd1407909, -25'd506847, -25'd2534237}, '{-25'd1464226, -25'd281582, 25'd2477921, -25'd619480, -25'd1351593}, '{25'd394215, 25'd1407909, 25'd3322666, 25'd619480, -25'd2759503}, '{25'd506847, 25'd450531, 25'd2590553, -25'd1407909, -25'd3435299}, '{-25'd1013695, 25'd337898, -25'd619480, -25'd1745808, -25'd2984768}}, '{'{-25'd1126328, -25'd506847, 25'd901062, -25'd1070011, -25'd844746}, '{-25'd1126328, -25'd1182644, -25'd281582, 25'd1126328, -25'd844746}, '{25'd281582, 25'd1238960, 25'd394215, -25'd1013695, -25'd619480}, '{-25'd394215, 25'd56316, 25'd619480, 25'd1238960, -25'd1013695}, '{-25'd1013695, 25'd1126328, -25'd1070011, -25'd450531, -25'd1126328}}, '{'{-25'd563164, 25'd168949, 25'd901062, 25'd732113, 25'd957378}, '{-25'd450531, 25'd1238960, 25'd168949, -25'd112633, -25'd225266}, '{25'd732113, 25'd901062, -25'd675797, -25'd56316, 25'd1070011}, '{-25'd1070011, 25'd112633, -25'd563164, 25'd506847, 25'd225266}, '{-25'd337898, 25'd281582, -25'd112633, -25'd337898, -25'd1013695}}, '{'{25'd957378, 25'd0, -25'd337898, 25'd1013695, -25'd1013695}, '{-25'd168949, 25'd0, 25'd1013695, 25'd168949, 25'd112633}, '{25'd1013695, 25'd56316, 25'd901062, -25'd1013695, 25'd788429}, '{-25'd394215, -25'd1126328, -25'd675797, 25'd1295277, 25'd844746}, '{25'd788429, 25'd901062, 25'd394215, 25'd957378, -25'd957378}}, '{'{25'd2703186, 25'd56316, -25'd1013695, -25'd1182644, 25'd0}, '{25'd1971073, -25'd1464226, -25'd2703186, -25'd957378, 25'd281582}, '{25'd337898, -25'd1464226, -25'd1802124, 25'd732113, 25'd1914757}, '{-25'd112633, -25'd1633175, -25'd1295277, 25'd563164, 25'd1914757}, '{25'd1126328, -25'd337898, -25'd506847, 25'd563164, 25'd1745808}}, '{'{-25'd844746, 25'd2703186, 25'd2646870, -25'd1182644, -25'd1182644}, '{-25'd168949, 25'd1858441, 25'd2534237, 25'd675797, -25'd281582}, '{25'd506847, 25'd2140022, 25'd4167412, 25'd450531, -25'd901062}, '{25'd1802124, 25'd1971073, 25'd4167412, 25'd1351593, 25'd1070011}, '{25'd732113, 25'd2534237, 25'd2308972, 25'd225266, -25'd675797}}, '{'{-25'd732113, -25'd506847, 25'd168949, 25'd225266, -25'd619480}, '{-25'd337898, 25'd788429, -25'd844746, 25'd394215, -25'd675797}, '{-25'd1858441, -25'd337898, -25'd168949, 25'd450531, 25'd225266}, '{-25'd1576859, -25'd732113, 25'd788429, 25'd112633, -25'd506847}, '{-25'd337898, -25'd563164, -25'd619480, 25'd225266, 25'd619480}}, '{'{-25'd563164, -25'd1070011, -25'd1182644, -25'd1126328, -25'd901062}, '{25'd788429, -25'd563164, -25'd450531, -25'd1182644, -25'd450531}, '{-25'd957378, -25'd337898, -25'd281582, -25'd1013695, -25'd56316}, '{-25'd394215, -25'd1126328, -25'd1013695, 25'd450531, -25'd844746}, '{25'd0, -25'd1182644, -25'd281582, 25'd957378, -25'd619480}}, '{'{-25'd506847, 25'd56316, 25'd619480, -25'd619480, 25'd619480}, '{-25'd112633, 25'd563164, 25'd619480, 25'd619480, 25'd56316}, '{25'd788429, 25'd732113, 25'd844746, 25'd619480, 25'd450531}, '{-25'd394215, -25'd168949, -25'd450531, -25'd168949, 25'd0}, '{25'd563164, -25'd506847, -25'd1238960, 25'd56316, 25'd281582}}, '{'{-25'd619480, -25'd563164, -25'd4280045, 25'd2703186, 25'd957378}, '{-25'd3153717, -25'd5293740, -25'd4786892, -25'd56316, -25'd1971073}, '{-25'd1689491, -25'd1182644, -25'd3773197, 25'd2477921, 25'd112633}, '{25'd337898, 25'd281582, -25'd844746, 25'd2759503, 25'd1013695}, '{25'd1126328, 25'd732113, -25'd1464226, 25'd3773197, 25'd3773197}}, '{'{25'd675797, 25'd2365288, 25'd732113, 25'd1126328, 25'd788429}, '{-25'd56316, 25'd225266, 25'd732113, 25'd1351593, 25'd225266}, '{-25'd1464226, -25'd1407909, 25'd394215, -25'd1013695, -25'd394215}, '{-25'd957378, 25'd450531, -25'd1295277, -25'd957378, -25'd394215}, '{25'd1126328, -25'd225266, -25'd337898, -25'd732113, 25'd788429}}, '{'{25'd675797, 25'd1351593, -25'd450531, 25'd394215, 25'd1576859}, '{-25'd337898, -25'd1070011, -25'd1745808, -25'd732113, -25'd56316}, '{25'd1576859, -25'd112633, -25'd394215, -25'd844746, -25'd56316}, '{25'd1126328, -25'd675797, -25'd1126328, 25'd1407909, -25'd788429}, '{25'd844746, -25'd788429, 25'd563164, 25'd1013695, 25'd1464226}}, '{'{-25'd225266, -25'd450531, 25'd901062, 25'd1351593, 25'd394215}, '{25'd506847, 25'd957378, -25'd1070011, -25'd901062, 25'd563164}, '{-25'd957378, -25'd56316, -25'd844746, -25'd844746, -25'd788429}, '{-25'd1070011, 25'd901062, 25'd901062, 25'd1013695, -25'd506847}, '{-25'd281582, -25'd1070011, -25'd394215, -25'd788429, 25'd337898}}, '{'{25'd281582, -25'd957378, -25'd1013695, 25'd0, 25'd901062}, '{25'd1182644, 25'd0, 25'd0, 25'd1070011, -25'd957378}, '{25'd1070011, 25'd563164, 25'd337898, 25'd337898, 25'd1238960}, '{25'd394215, -25'd394215, 25'd1013695, 25'd225266, 25'd619480}, '{25'd450531, -25'd56316, 25'd844746, -25'd394215, -25'd394215}}, '{'{-25'd225266, -25'd337898, 25'd225266, -25'd168949, -25'd56316}, '{25'd732113, 25'd1238960, -25'd1126328, 25'd901062, -25'd1126328}, '{25'd281582, 25'd337898, -25'd225266, -25'd112633, -25'd394215}, '{-25'd394215, 25'd0, -25'd1295277, -25'd281582, -25'd506847}, '{-25'd225266, 25'd1182644, 25'd1126328, 25'd1295277, 25'd1070011}}, '{'{-25'd168949, -25'd1070011, 25'd2928452, 25'd4617943, -25'd1126328}, '{25'd619480, 25'd450531, 25'd3266350, 25'd4167412, 25'd0}, '{-25'd1464226, -25'd1858441, 25'd2308972, 25'd4448994, -25'd2534237}, '{-25'd1351593, -25'd2308972, 25'd1070011, 25'd2984768, -25'd2196339}, '{-25'd2815819, -25'd3435299, -25'd732113, -25'd225266, -25'd5124791}}, '{'{-25'd1802124, -25'd56316, 25'd1576859, -25'd1802124, -25'd1633175}, '{-25'd225266, 25'd0, 25'd2646870, -25'd281582, -25'd619480}, '{25'd901062, 25'd1633175, 25'd2984768, 25'd2590553, 25'd1407909}, '{25'd1745808, 25'd2027390, 25'd1971073, 25'd2646870, 25'd0}, '{25'd1013695, 25'd2534237, 25'd1914757, 25'd2083706, 25'd732113}}, '{'{-25'd957378, 25'd1013695, 25'd788429, 25'd619480, 25'd225266}, '{-25'd1126328, -25'd1070011, -25'd732113, 25'd675797, 25'd506847}, '{25'd1013695, 25'd394215, 25'd1182644, 25'd844746, 25'd168949}, '{25'd0, 25'd1182644, -25'd901062, -25'd1070011, -25'd112633}, '{25'd450531, 25'd56316, -25'd1013695, 25'd1295277, 25'd1126328}}, '{'{25'd337898, -25'd168949, 25'd168949, 25'd563164, 25'd450531}, '{25'd732113, 25'd563164, 25'd732113, 25'd1126328, -25'd1182644}, '{-25'd506847, 25'd450531, 25'd1576859, 25'd1633175, -25'd1464226}, '{-25'd112633, 25'd281582, 25'd732113, 25'd506847, -25'd394215}, '{-25'd168949, 25'd1126328, 25'd1351593, 25'd281582, 25'd506847}}, '{'{-25'd675797, 25'd112633, 25'd337898, -25'd1070011, 25'd281582}, '{-25'd1126328, 25'd1238960, -25'd675797, -25'd506847, 25'd788429}, '{-25'd1126328, 25'd1013695, -25'd788429, -25'd1013695, 25'd1013695}, '{25'd1013695, -25'd844746, -25'd450531, -25'd1070011, 25'd675797}, '{25'd1182644, 25'd788429, -25'd901062, -25'd1182644, -25'd1070011}}, '{'{25'd675797, -25'd563164, 25'd450531, 25'd788429, -25'd56316}, '{-25'd168949, -25'd1126328, 25'd450531, -25'd112633, 25'd225266}, '{25'd1070011, 25'd844746, 25'd844746, -25'd1013695, 25'd1182644}, '{25'd450531, -25'd506847, 25'd1238960, -25'd788429, -25'd1295277}, '{-25'd337898, -25'd168949, -25'd844746, 25'd1013695, 25'd1126328}}, '{'{25'd56316, -25'd563164, -25'd394215, 25'd1295277, 25'd281582}, '{-25'd957378, 25'd619480, 25'd1013695, 25'd168949, 25'd337898}, '{25'd675797, 25'd168949, 25'd563164, -25'd1126328, 25'd675797}, '{25'd1126328, -25'd1013695, 25'd225266, -25'd1126328, 25'd337898}, '{-25'd225266, 25'd112633, 25'd563164, 25'd1238960, -25'd56316}}, '{'{-25'd394215, 25'd563164, 25'd1407909, 25'd1520542, 25'd168949}, '{25'd112633, -25'd337898, 25'd957378, 25'd1914757, 25'd1407909}, '{25'd1013695, 25'd2027390, 25'd1070011, 25'd168949, 25'd1520542}, '{25'd732113, 25'd563164, 25'd732113, -25'd1182644, -25'd788429}, '{25'd1238960, -25'd56316, 25'd450531, 25'd563164, 25'd563164}}, '{'{25'd56316, 25'd1576859, 25'd563164, 25'd2477921, -25'd6251118}, '{25'd844746, 25'd1013695, 25'd2872135, 25'd4336361, 25'd1013695}, '{25'd2140022, 25'd675797, 25'd1576859, 25'd2534237, 25'd1126328}, '{25'd112633, -25'd1971073, -25'd394215, 25'd844746, 25'd0}, '{25'd56316, 25'd450531, -25'd2252655, 25'd394215, -25'd281582}}, '{'{-25'd675797, -25'd1126328, -25'd675797, 25'd0, -25'd112633}, '{25'd281582, -25'd337898, 25'd1013695, 25'd450531, 25'd1182644}, '{25'd2815819, 25'd2027390, 25'd2815819, 25'd3435299, 25'd675797}, '{25'd1914757, 25'd2703186, 25'd3435299, 25'd2646870, -25'd1633175}, '{25'd1633175, 25'd1351593, 25'd1914757, -25'd1802124, -25'd7208497}}}
};
