localparam bit signed [0:10][15:0] Output3 = '{16'd21523, 16'd25074, -16'd11610, -16'd29433, 16'd6102, -16'd17479, 16'd27563, -16'd936, 16'd5069, 16'd17281, 16'd32478};
