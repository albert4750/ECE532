localparam bit signed [0:31][0:63][0:0][0:0][24:0] Weight2 = '{
    '{'{'{25'd581}}, '{'{-25'd3873}}, '{'{-25'd1033}}, '{'{-25'd8197}}, '{'{25'd194}}, '{'{25'd1355}}, '{'{-25'd1485}}, '{'{25'd1807}}, '{'{25'd1355}}, '{'{-25'd2582}}, '{'{-25'd3356}}, '{'{-25'd1291}}, '{'{-25'd2195}}, '{'{25'd1936}}, '{'{-25'd3808}}, '{'{25'd1226}}, '{'{-25'd65}}, '{'{-25'd4389}}, '{'{-25'd3615}}, '{'{25'd452}}, '{'{-25'd2130}}, '{'{25'd904}}, '{'{25'd3744}}, '{'{-25'd2453}}, '{'{-25'd1097}}, '{'{25'd3486}}, '{'{-25'd904}}, '{'{25'd4776}}, '{'{25'd4325}}, '{'{25'd2324}}, '{'{-25'd1807}}, '{'{-25'd387}}, '{'{-25'd1549}}, '{'{-25'd5551}}, '{'{25'd1614}}, '{'{-25'd129}}, '{'{-25'd4325}}, '{'{25'd839}}, '{'{-25'd3421}}, '{'{-25'd5551}}, '{'{25'd1872}}, '{'{-25'd323}}, '{'{-25'd5680}}, '{'{25'd4583}}, '{'{-25'd1033}}, '{'{25'd2969}}, '{'{25'd1872}}, '{'{-25'd2646}}, '{'{-25'd3421}}, '{'{-25'd3486}}, '{'{25'd0}}, '{'{25'd4906}}, '{'{-25'd1743}}, '{'{25'd387}}, '{'{-25'd387}}, '{'{25'd1743}}, '{'{25'd1226}}, '{'{25'd0}}, '{'{25'd1291}}, '{'{-25'd5035}}, '{'{-25'd2453}}, '{'{-25'd3744}}, '{'{-25'd2066}}, '{'{-25'd2711}}},
    '{'{'{-25'd3761}}, '{'{-25'd3352}}, '{'{-25'd7440}}, '{'{-25'd9238}}, '{'{-25'd10301}}, '{'{25'd1226}}, '{'{-25'd3188}}, '{'{-25'd3842}}, '{'{-25'd1635}}, '{'{-25'd82}}, '{'{-25'd4170}}, '{'{25'd1553}}, '{'{-25'd1145}}, '{'{25'd4088}}, '{'{25'd1553}}, '{'{25'd2616}}, '{'{25'd5478}}, '{'{-25'd5559}}, '{'{-25'd245}}, '{'{-25'd2780}}, '{'{-25'd1717}}, '{'{25'd4415}}, '{'{-25'd3842}}, '{'{-25'd82}}, '{'{25'd4415}}, '{'{-25'd2780}}, '{'{25'd164}}, '{'{25'd1390}}, '{'{25'd3270}}, '{'{-25'd4006}}, '{'{25'd4415}}, '{'{-25'd1635}}, '{'{25'd5232}}, '{'{25'd2616}}, '{'{-25'd3597}}, '{'{-25'd8421}}, '{'{25'd5232}}, '{'{25'd1553}}, '{'{25'd4006}}, '{'{-25'd9647}}, '{'{-25'd2371}}, '{'{25'd10383}}, '{'{25'd3352}}, '{'{25'd4660}}, '{'{25'd2044}}, '{'{25'd4905}}, '{'{-25'd2289}}, '{'{25'd5886}}, '{'{-25'd4170}}, '{'{25'd899}}, '{'{25'd2780}}, '{'{-25'd1145}}, '{'{-25'd4824}}, '{'{-25'd2616}}, '{'{-25'd3025}}, '{'{25'd0}}, '{'{25'd2453}}, '{'{25'd2616}}, '{'{-25'd2126}}, '{'{-25'd3515}}, '{'{25'd10056}}, '{'{-25'd1635}}, '{'{25'd4905}}, '{'{-25'd4333}}},
    '{'{'{25'd6546}}, '{'{25'd1021}}, '{'{-25'd1561}}, '{'{25'd6125}}, '{'{-25'd1922}}, '{'{25'd2943}}, '{'{25'd5525}}, '{'{-25'd540}}, '{'{25'd1741}}, '{'{-25'd7566}}, '{'{25'd1441}}, '{'{-25'd3663}}, '{'{-25'd2943}}, '{'{-25'd2162}}, '{'{25'd4864}}, '{'{-25'd1021}}, '{'{25'd3783}}, '{'{-25'd5044}}, '{'{25'd1141}}, '{'{-25'd1561}}, '{'{-25'd120}}, '{'{-25'd300}}, '{'{-25'd3543}}, '{'{-25'd1321}}, '{'{25'd2882}}, '{'{-25'd2822}}, '{'{-25'd2762}}, '{'{25'd3183}}, '{'{25'd4264}}, '{'{-25'd240}}, '{'{25'd3003}}, '{'{25'd3963}}, '{'{-25'd3423}}, '{'{-25'd5525}}, '{'{-25'd901}}, '{'{-25'd1802}}, '{'{-25'd2162}}, '{'{25'd240}}, '{'{-25'd3303}}, '{'{-25'd7687}}, '{'{-25'd3543}}, '{'{25'd4624}}, '{'{25'd1741}}, '{'{-25'd3123}}, '{'{-25'd2522}}, '{'{25'd3723}}, '{'{25'd1321}}, '{'{25'd3123}}, '{'{25'd2042}}, '{'{-25'd4804}}, '{'{-25'd3903}}, '{'{25'd1501}}, '{'{-25'd1441}}, '{'{25'd2822}}, '{'{-25'd1681}}, '{'{-25'd2042}}, '{'{-25'd1922}}, '{'{-25'd2042}}, '{'{25'd4864}}, '{'{-25'd4444}}, '{'{25'd0}}, '{'{-25'd901}}, '{'{25'd2462}}, '{'{25'd4744}}},
    '{'{'{25'd3394}}, '{'{-25'd1048}}, '{'{-25'd2845}}, '{'{-25'd599}}, '{'{25'd1098}}, '{'{25'd2745}}, '{'{-25'd3045}}, '{'{-25'd2596}}, '{'{25'd399}}, '{'{25'd6239}}, '{'{-25'd749}}, '{'{25'd250}}, '{'{-25'd1697}}, '{'{-25'd2945}}, '{'{25'd5391}}, '{'{-25'd3195}}, '{'{25'd3843}}, '{'{-25'd4692}}, '{'{-25'd4842}}, '{'{25'd3893}}, '{'{25'd2196}}, '{'{-25'd4792}}, '{'{-25'd2945}}, '{'{25'd6289}}, '{'{25'd3195}}, '{'{25'd799}}, '{'{-25'd1148}}, '{'{25'd2396}}, '{'{25'd1348}}, '{'{25'd1497}}, '{'{-25'd2645}}, '{'{-25'd499}}, '{'{-25'd3494}}, '{'{-25'd1298}}, '{'{-25'd5041}}, '{'{25'd4642}}, '{'{-25'd6339}}, '{'{25'd50}}, '{'{25'd3145}}, '{'{-25'd3145}}, '{'{25'd2745}}, '{'{-25'd5241}}, '{'{-25'd948}}, '{'{-25'd2396}}, '{'{-25'd4892}}, '{'{25'd1198}}, '{'{25'd4243}}, '{'{25'd2396}}, '{'{-25'd3494}}, '{'{-25'd5690}}, '{'{25'd2895}}, '{'{25'd2695}}, '{'{25'd1398}}, '{'{-25'd2096}}, '{'{-25'd6389}}, '{'{25'd3943}}, '{'{-25'd4243}}, '{'{25'd449}}, '{'{25'd1647}}, '{'{-25'd299}}, '{'{25'd2496}}, '{'{25'd200}}, '{'{25'd699}}, '{'{25'd3644}}},
    '{'{'{25'd8638}}, '{'{25'd1212}}, '{'{-25'd303}}, '{'{25'd6971}}, '{'{25'd1970}}, '{'{25'd303}}, '{'{-25'd455}}, '{'{-25'd1061}}, '{'{-25'd2273}}, '{'{25'd8638}}, '{'{-25'd8183}}, '{'{25'd1061}}, '{'{-25'd303}}, '{'{-25'd1818}}, '{'{25'd5910}}, '{'{-25'd4698}}, '{'{25'd19246}}, '{'{25'd5304}}, '{'{-25'd3334}}, '{'{25'd6213}}, '{'{25'd1818}}, '{'{25'd758}}, '{'{-25'd3940}}, '{'{-25'd6516}}, '{'{25'd3637}}, '{'{25'd1364}}, '{'{25'd3182}}, '{'{-25'd2425}}, '{'{-25'd2425}}, '{'{25'd3637}}, '{'{-25'd2576}}, '{'{25'd2425}}, '{'{-25'd4092}}, '{'{25'd303}}, '{'{-25'd3940}}, '{'{-25'd2273}}, '{'{25'd2425}}, '{'{25'd5304}}, '{'{-25'd3485}}, '{'{-25'd5304}}, '{'{-25'd5152}}, '{'{25'd14093}}, '{'{-25'd2879}}, '{'{-25'd758}}, '{'{25'd3182}}, '{'{-25'd3637}}, '{'{25'd1364}}, '{'{25'd4395}}, '{'{25'd909}}, '{'{-25'd3182}}, '{'{-25'd3485}}, '{'{-25'd4092}}, '{'{25'd1364}}, '{'{-25'd3334}}, '{'{-25'd3940}}, '{'{25'd1061}}, '{'{-25'd5304}}, '{'{25'd3485}}, '{'{-25'd1818}}, '{'{25'd2728}}, '{'{-25'd1818}}, '{'{25'd4395}}, '{'{25'd0}}, '{'{-25'd1970}}},
    '{'{'{25'd2316}}, '{'{25'd2920}}, '{'{-25'd805}}, '{'{25'd604}}, '{'{-25'd2819}}, '{'{25'd0}}, '{'{-25'd1913}}, '{'{25'd9162}}, '{'{-25'd101}}, '{'{-25'd1007}}, '{'{25'd101}}, '{'{-25'd4128}}, '{'{-25'd4933}}, '{'{25'd302}}, '{'{25'd2920}}, '{'{25'd403}}, '{'{25'd302}}, '{'{-25'd2618}}, '{'{-25'd6544}}, '{'{25'd1208}}, '{'{-25'd4228}}, '{'{25'd2718}}, '{'{25'd2618}}, '{'{-25'd3725}}, '{'{25'd5135}}, '{'{-25'd3020}}, '{'{25'd4732}}, '{'{-25'd6141}}, '{'{-25'd5336}}, '{'{25'd7551}}, '{'{-25'd2114}}, '{'{-25'd2114}}, '{'{-25'd201}}, '{'{25'd1409}}, '{'{25'd4027}}, '{'{25'd2316}}, '{'{25'd5437}}, '{'{25'd0}}, '{'{-25'd3524}}, '{'{25'd4732}}, '{'{25'd3322}}, '{'{25'd12786}}, '{'{25'd705}}, '{'{-25'd1007}}, '{'{-25'd4631}}, '{'{-25'd4128}}, '{'{-25'd302}}, '{'{25'd6343}}, '{'{-25'd7148}}, '{'{-25'd3725}}, '{'{-25'd3121}}, '{'{-25'd6947}}, '{'{25'd1611}}, '{'{-25'd1812}}, '{'{-25'd1611}}, '{'{-25'd8457}}, '{'{25'd906}}, '{'{25'd7148}}, '{'{-25'd6947}}, '{'{25'd4228}}, '{'{-25'd1107}}, '{'{25'd6242}}, '{'{-25'd2517}}, '{'{25'd3121}}},
    '{'{'{-25'd2903}}, '{'{25'd0}}, '{'{25'd2516}}, '{'{-25'd8259}}, '{'{25'd903}}, '{'{-25'd903}}, '{'{25'd4452}}, '{'{25'd5807}}, '{'{25'd4323}}, '{'{-25'd4645}}, '{'{-25'd6646}}, '{'{-25'd839}}, '{'{-25'd194}}, '{'{-25'd1290}}, '{'{25'd4129}}, '{'{25'd4323}}, '{'{25'd2839}}, '{'{25'd4968}}, '{'{25'd3549}}, '{'{25'd1936}}, '{'{25'd5033}}, '{'{-25'd2774}}, '{'{-25'd1097}}, '{'{-25'd2839}}, '{'{25'd2000}}, '{'{25'd3807}}, '{'{25'd3549}}, '{'{-25'd3678}}, '{'{-25'd4581}}, '{'{25'd4129}}, '{'{25'd2774}}, '{'{25'd5162}}, '{'{25'd5420}}, '{'{-25'd2839}}, '{'{-25'd4194}}, '{'{25'd1613}}, '{'{-25'd4387}}, '{'{25'd1097}}, '{'{25'd2903}}, '{'{-25'd6323}}, '{'{-25'd2323}}, '{'{25'd4775}}, '{'{-25'd4258}}, '{'{-25'd1419}}, '{'{25'd2452}}, '{'{25'd258}}, '{'{25'd3678}}, '{'{25'd8065}}, '{'{-25'd903}}, '{'{25'd516}}, '{'{25'd323}}, '{'{-25'd839}}, '{'{-25'd3742}}, '{'{25'd1548}}, '{'{-25'd5033}}, '{'{25'd1419}}, '{'{25'd5226}}, '{'{-25'd2516}}, '{'{25'd1161}}, '{'{-25'd4323}}, '{'{25'd2387}}, '{'{25'd6258}}, '{'{25'd2710}}, '{'{25'd2452}}},
    '{'{'{-25'd2241}}, '{'{25'd1027}}, '{'{25'd2708}}, '{'{25'd1214}}, '{'{25'd3082}}, '{'{-25'd747}}, '{'{25'd3175}}, '{'{-25'd5136}}, '{'{25'd467}}, '{'{25'd7004}}, '{'{25'd1401}}, '{'{25'd1681}}, '{'{-25'd2708}}, '{'{-25'd1121}}, '{'{25'd5323}}, '{'{-25'd3829}}, '{'{-25'd4950}}, '{'{25'd1214}}, '{'{25'd3082}}, '{'{25'd3829}}, '{'{25'd4669}}, '{'{25'd2055}}, '{'{-25'd560}}, '{'{25'd374}}, '{'{-25'd4202}}, '{'{-25'd3922}}, '{'{25'd3269}}, '{'{-25'd2708}}, '{'{-25'd2521}}, '{'{-25'd654}}, '{'{25'd4576}}, '{'{-25'd2708}}, '{'{25'd1681}}, '{'{25'd1401}}, '{'{25'd4109}}, '{'{-25'd1307}}, '{'{25'd3549}}, '{'{25'd4763}}, '{'{-25'd3269}}, '{'{25'd3922}}, '{'{25'd560}}, '{'{-25'd1588}}, '{'{-25'd1214}}, '{'{25'd2521}}, '{'{25'd560}}, '{'{-25'd1121}}, '{'{-25'd187}}, '{'{-25'd2055}}, '{'{25'd93}}, '{'{25'd11860}}, '{'{-25'd5136}}, '{'{25'd1494}}, '{'{25'd4296}}, '{'{25'd1027}}, '{'{-25'd3642}}, '{'{-25'd2055}}, '{'{-25'd2708}}, '{'{-25'd5883}}, '{'{25'd3455}}, '{'{-25'd187}}, '{'{25'd3736}}, '{'{25'd2895}}, '{'{-25'd467}}, '{'{25'd2148}}},
    '{'{'{25'd6132}}, '{'{-25'd6059}}, '{'{25'd0}}, '{'{-25'd9344}}, '{'{25'd73}}, '{'{25'd5110}}, '{'{25'd4161}}, '{'{25'd219}}, '{'{25'd4964}}, '{'{-25'd2701}}, '{'{25'd2774}}, '{'{-25'd2774}}, '{'{-25'd2336}}, '{'{25'd1460}}, '{'{-25'd3650}}, '{'{-25'd1168}}, '{'{25'd6497}}, '{'{-25'd4453}}, '{'{25'd3066}}, '{'{25'd5256}}, '{'{25'd73}}, '{'{25'd2336}}, '{'{-25'd1387}}, '{'{25'd657}}, '{'{-25'd5037}}, '{'{25'd3869}}, '{'{25'd4599}}, '{'{25'd1533}}, '{'{-25'd2044}}, '{'{25'd2190}}, '{'{25'd2847}}, '{'{25'd3066}}, '{'{25'd1460}}, '{'{-25'd4964}}, '{'{25'd2409}}, '{'{-25'd3796}}, '{'{-25'd3066}}, '{'{25'd73}}, '{'{25'd5548}}, '{'{-25'd7519}}, '{'{-25'd2336}}, '{'{25'd3796}}, '{'{25'd3139}}, '{'{-25'd1971}}, '{'{25'd1533}}, '{'{25'd3212}}, '{'{-25'd511}}, '{'{25'd2117}}, '{'{25'd4088}}, '{'{-25'd1533}}, '{'{-25'd219}}, '{'{-25'd2628}}, '{'{25'd5548}}, '{'{-25'd2190}}, '{'{25'd2044}}, '{'{-25'd1314}}, '{'{25'd4380}}, '{'{-25'd1679}}, '{'{-25'd3066}}, '{'{25'd3212}}, '{'{-25'd1606}}, '{'{-25'd803}}, '{'{-25'd511}}, '{'{25'd4526}}},
    '{'{'{25'd996}}, '{'{-25'd5103}}, '{'{-25'd2116}}, '{'{25'd311}}, '{'{-25'd7903}}, '{'{25'd4979}}, '{'{25'd6223}}, '{'{25'd4481}}, '{'{25'd5788}}, '{'{25'd1991}}, '{'{25'd1120}}, '{'{25'd1556}}, '{'{-25'd933}}, '{'{25'd996}}, '{'{25'd3423}}, '{'{25'd6846}}, '{'{25'd747}}, '{'{-25'd1120}}, '{'{25'd1618}}, '{'{25'd5227}}, '{'{25'd809}}, '{'{25'd560}}, '{'{25'd4170}}, '{'{-25'd4418}}, '{'{-25'd3547}}, '{'{-25'd1680}}, '{'{-25'd6099}}, '{'{-25'd560}}, '{'{-25'd311}}, '{'{-25'd4916}}, '{'{-25'd3112}}, '{'{25'd373}}, '{'{-25'd4730}}, '{'{-25'd4854}}, '{'{-25'd1369}}, '{'{25'd2925}}, '{'{-25'd1618}}, '{'{-25'd1556}}, '{'{-25'd2427}}, '{'{-25'd7468}}, '{'{25'd1618}}, '{'{-25'd3983}}, '{'{25'd1556}}, '{'{-25'd4107}}, '{'{25'd5476}}, '{'{-25'd187}}, '{'{-25'd2178}}, '{'{25'd4107}}, '{'{-25'd933}}, '{'{25'd2178}}, '{'{-25'd2116}}, '{'{-25'd5663}}, '{'{25'd5290}}, '{'{-25'd933}}, '{'{-25'd1120}}, '{'{25'd1805}}, '{'{-25'd3921}}, '{'{-25'd5103}}, '{'{-25'd1245}}, '{'{25'd3423}}, '{'{25'd1307}}, '{'{-25'd2303}}, '{'{-25'd2676}}, '{'{25'd124}}},
    '{'{'{25'd1034}}, '{'{-25'd969}}, '{'{-25'd6720}}, '{'{-25'd8271}}, '{'{25'd3554}}, '{'{25'd4071}}, '{'{25'd4976}}, '{'{25'd5622}}, '{'{-25'd452}}, '{'{-25'd1809}}, '{'{-25'd5363}}, '{'{-25'd2585}}, '{'{-25'd1939}}, '{'{25'd3296}}, '{'{-25'd3166}}, '{'{-25'd129}}, '{'{25'd5105}}, '{'{25'd1809}}, '{'{25'd2585}}, '{'{25'd3683}}, '{'{25'd3360}}, '{'{-25'd2908}}, '{'{25'd1292}}, '{'{-25'd4459}}, '{'{-25'd1292}}, '{'{-25'd4976}}, '{'{-25'd2132}}, '{'{-25'd2779}}, '{'{25'd4911}}, '{'{25'd1551}}, '{'{25'd5170}}, '{'{25'd4911}}, '{'{25'd3166}}, '{'{25'd969}}, '{'{-25'd7431}}, '{'{-25'd6914}}, '{'{-25'd194}}, '{'{-25'd3425}}, '{'{25'd1163}}, '{'{25'd646}}, '{'{-25'd4006}}, '{'{25'd3296}}, '{'{25'd1486}}, '{'{-25'd2003}}, '{'{25'd5170}}, '{'{-25'd4523}}, '{'{-25'd2326}}, '{'{25'd3748}}, '{'{-25'd1809}}, '{'{-25'd1680}}, '{'{25'd452}}, '{'{-25'd1357}}, '{'{-25'd3296}}, '{'{-25'd5040}}, '{'{-25'd5557}}, '{'{-25'd1874}}, '{'{25'd2456}}, '{'{-25'd194}}, '{'{-25'd1680}}, '{'{25'd1874}}, '{'{-25'd840}}, '{'{-25'd2132}}, '{'{25'd4847}}, '{'{-25'd4330}}},
    '{'{'{25'd1980}}, '{'{25'd888}}, '{'{25'd2048}}, '{'{-25'd410}}, '{'{25'd683}}, '{'{25'd1570}}, '{'{25'd4643}}, '{'{25'd1229}}, '{'{-25'd4506}}, '{'{-25'd7784}}, '{'{-25'd6623}}, '{'{-25'd2253}}, '{'{25'd4438}}, '{'{-25'd341}}, '{'{-25'd205}}, '{'{-25'd1844}}, '{'{25'd5940}}, '{'{25'd3141}}, '{'{25'd2731}}, '{'{-25'd3550}}, '{'{-25'd3004}}, '{'{25'd2731}}, '{'{25'd478}}, '{'{-25'd4302}}, '{'{-25'd1502}}, '{'{25'd2595}}, '{'{25'd2390}}, '{'{-25'd273}}, '{'{-25'd683}}, '{'{25'd3619}}, '{'{25'd3209}}, '{'{-25'd205}}, '{'{-25'd1434}}, '{'{25'd2868}}, '{'{25'd2526}}, '{'{-25'd2117}}, '{'{-25'd4302}}, '{'{-25'd1570}}, '{'{25'd2321}}, '{'{-25'd8740}}, '{'{-25'd3004}}, '{'{25'd7579}}, '{'{-25'd888}}, '{'{-25'd1502}}, '{'{-25'd1297}}, '{'{25'd3277}}, '{'{25'd4097}}, '{'{-25'd4643}}, '{'{25'd1570}}, '{'{-25'd2526}}, '{'{25'd3619}}, '{'{-25'd3141}}, '{'{-25'd4370}}, '{'{-25'd1502}}, '{'{-25'd4916}}, '{'{-25'd3073}}, '{'{-25'd1775}}, '{'{25'd6760}}, '{'{25'd3687}}, '{'{25'd341}}, '{'{-25'd2321}}, '{'{-25'd546}}, '{'{-25'd4506}}, '{'{25'd3073}}},
    '{'{'{25'd7837}}, '{'{-25'd2689}}, '{'{-25'd3381}}, '{'{25'd1614}}, '{'{25'd6454}}, '{'{25'd4226}}, '{'{-25'd2459}}, '{'{-25'd538}}, '{'{25'd307}}, '{'{-25'd1383}}, '{'{-25'd7607}}, '{'{-25'd2612}}, '{'{25'd1614}}, '{'{-25'd5302}}, '{'{25'd6531}}, '{'{-25'd2997}}, '{'{25'd9758}}, '{'{25'd4226}}, '{'{25'd3227}}, '{'{-25'd2920}}, '{'{25'd1998}}, '{'{25'd4380}}, '{'{-25'd3765}}, '{'{25'd6992}}, '{'{-25'd5532}}, '{'{-25'd1767}}, '{'{-25'd1460}}, '{'{-25'd4380}}, '{'{25'd1153}}, '{'{-25'd1921}}, '{'{25'd692}}, '{'{-25'd4917}}, '{'{-25'd2689}}, '{'{25'd2843}}, '{'{-25'd1844}}, '{'{-25'd1767}}, '{'{25'd3304}}, '{'{25'd768}}, '{'{25'd538}}, '{'{-25'd6224}}, '{'{-25'd9681}}, '{'{25'd5532}}, '{'{-25'd1690}}, '{'{-25'd8682}}, '{'{-25'd3073}}, '{'{-25'd692}}, '{'{25'd3304}}, '{'{25'd2766}}, '{'{25'd2151}}, '{'{-25'd1306}}, '{'{25'd4226}}, '{'{-25'd922}}, '{'{25'd4841}}, '{'{25'd4303}}, '{'{25'd3227}}, '{'{25'd1998}}, '{'{25'd4610}}, '{'{25'd8913}}, '{'{-25'd3611}}, '{'{-25'd2382}}, '{'{-25'd154}}, '{'{-25'd768}}, '{'{-25'd2305}}, '{'{25'd3765}}},
    '{'{'{25'd5904}}, '{'{25'd293}}, '{'{25'd4440}}, '{'{25'd1122}}, '{'{25'd4587}}, '{'{25'd5270}}, '{'{25'd98}}, '{'{25'd1025}}, '{'{-25'd488}}, '{'{-25'd4343}}, '{'{-25'd2293}}, '{'{-25'd4489}}, '{'{-25'd1122}}, '{'{-25'd2976}}, '{'{-25'd1952}}, '{'{-25'd195}}, '{'{25'd6197}}, '{'{25'd2635}}, '{'{-25'd2391}}, '{'{25'd2293}}, '{'{25'd2830}}, '{'{25'd4147}}, '{'{25'd537}}, '{'{-25'd4831}}, '{'{25'd2928}}, '{'{25'd586}}, '{'{25'd3269}}, '{'{25'd1757}}, '{'{25'd3757}}, '{'{25'd2537}}, '{'{25'd4928}}, '{'{25'd146}}, '{'{-25'd3904}}, '{'{-25'd2586}}, '{'{-25'd1171}}, '{'{25'd4147}}, '{'{25'd2976}}, '{'{25'd4440}}, '{'{-25'd488}}, '{'{-25'd6050}}, '{'{-25'd3220}}, '{'{25'd5953}}, '{'{-25'd5563}}, '{'{25'd2245}}, '{'{-25'd1025}}, '{'{25'd3269}}, '{'{25'd4684}}, '{'{25'd2098}}, '{'{25'd293}}, '{'{-25'd6099}}, '{'{-25'd1171}}, '{'{25'd3123}}, '{'{-25'd3416}}, '{'{-25'd878}}, '{'{25'd2049}}, '{'{-25'd2147}}, '{'{-25'd1610}}, '{'{25'd2879}}, '{'{25'd3074}}, '{'{-25'd3367}}, '{'{-25'd1122}}, '{'{-25'd2537}}, '{'{25'd3952}}, '{'{-25'd634}}},
    '{'{'{25'd3436}}, '{'{-25'd1826}}, '{'{-25'd3544}}, '{'{-25'd1772}}, '{'{-25'd322}}, '{'{25'd1181}}, '{'{-25'd4134}}, '{'{25'd2416}}, '{'{-25'd1664}}, '{'{-25'd805}}, '{'{-25'd3651}}, '{'{25'd3759}}, '{'{25'd5316}}, '{'{25'd3759}}, '{'{25'd4134}}, '{'{25'd4510}}, '{'{25'd4564}}, '{'{-25'd3329}}, '{'{25'd4295}}, '{'{25'd859}}, '{'{-25'd1826}}, '{'{25'd1772}}, '{'{25'd2470}}, '{'{-25'd6228}}, '{'{25'd2470}}, '{'{25'd4940}}, '{'{-25'd5853}}, '{'{25'd1074}}, '{'{-25'd913}}, '{'{25'd5369}}, '{'{-25'd4081}}, '{'{25'd4403}}, '{'{25'd3329}}, '{'{25'd2255}}, '{'{-25'd483}}, '{'{-25'd4779}}, '{'{-25'd2255}}, '{'{25'd5208}}, '{'{-25'd3007}}, '{'{-25'd3866}}, '{'{-25'd2255}}, '{'{25'd2201}}, '{'{25'd1235}}, '{'{-25'd537}}, '{'{25'd4403}}, '{'{-25'd3007}}, '{'{-25'd5262}}, '{'{-25'd805}}, '{'{-25'd2309}}, '{'{-25'd6873}}, '{'{-25'd4510}}, '{'{-25'd1074}}, '{'{25'd1879}}, '{'{25'd2362}}, '{'{25'd644}}, '{'{25'd2201}}, '{'{25'd2792}}, '{'{25'd4027}}, '{'{-25'd3973}}, '{'{25'd805}}, '{'{25'd3544}}, '{'{25'd2631}}, '{'{25'd3651}}, '{'{-25'd4618}}},
    '{'{'{-25'd8729}}, '{'{25'd0}}, '{'{25'd153}}, '{'{25'd613}}, '{'{25'd12863}}, '{'{-25'd2450}}, '{'{-25'd1838}}, '{'{-25'd1072}}, '{'{-25'd3063}}, '{'{-25'd2603}}, '{'{-25'd4135}}, '{'{-25'd4441}}, '{'{25'd5666}}, '{'{25'd6585}}, '{'{25'd4594}}, '{'{-25'd13782}}, '{'{25'd1378}}, '{'{-25'd2910}}, '{'{25'd613}}, '{'{-25'd459}}, '{'{-25'd3522}}, '{'{-25'd5207}}, '{'{-25'd7504}}, '{'{25'd3675}}, '{'{25'd15313}}, '{'{25'd1072}}, '{'{-25'd2144}}, '{'{25'd5207}}, '{'{-25'd2297}}, '{'{25'd0}}, '{'{-25'd4441}}, '{'{25'd3369}}, '{'{25'd2603}}, '{'{25'd16232}}, '{'{-25'd766}}, '{'{25'd7504}}, '{'{25'd5513}}, '{'{25'd613}}, '{'{25'd2297}}, '{'{25'd0}}, '{'{25'd3369}}, '{'{25'd6585}}, '{'{-25'd1225}}, '{'{-25'd3982}}, '{'{-25'd3982}}, '{'{-25'd4441}}, '{'{-25'd5666}}, '{'{-25'd9341}}, '{'{25'd5819}}, '{'{-25'd3216}}, '{'{-25'd3675}}, '{'{-25'd459}}, '{'{-25'd613}}, '{'{-25'd3522}}, '{'{-25'd7197}}, '{'{25'd5972}}, '{'{-25'd5053}}, '{'{25'd19448}}, '{'{-25'd2910}}, '{'{25'd4594}}, '{'{25'd4135}}, '{'{25'd459}}, '{'{25'd1225}}, '{'{-25'd2297}}},
    '{'{'{25'd6928}}, '{'{25'd4730}}, '{'{25'd600}}, '{'{-25'd7395}}, '{'{-25'd7195}}, '{'{-25'd999}}, '{'{25'd3931}}, '{'{25'd3797}}, '{'{25'd933}}, '{'{25'd200}}, '{'{25'd3931}}, '{'{-25'd6795}}, '{'{-25'd4330}}, '{'{25'd666}}, '{'{-25'd2998}}, '{'{-25'd3597}}, '{'{-25'd2532}}, '{'{25'd2865}}, '{'{-25'd4663}}, '{'{25'd2398}}, '{'{-25'd799}}, '{'{-25'd4197}}, '{'{25'd7728}}, '{'{-25'd933}}, '{'{25'd600}}, '{'{-25'd2198}}, '{'{-25'd6862}}, '{'{25'd1266}}, '{'{-25'd6662}}, '{'{25'd2265}}, '{'{-25'd666}}, '{'{-25'd133}}, '{'{25'd3131}}, '{'{-25'd8527}}, '{'{25'd799}}, '{'{-25'd2998}}, '{'{-25'd4597}}, '{'{25'd1799}}, '{'{-25'd4930}}, '{'{-25'd1732}}, '{'{25'd1932}}, '{'{-25'd8527}}, '{'{-25'd1332}}, '{'{25'd5729}}, '{'{-25'd1332}}, '{'{-25'd2931}}, '{'{-25'd2332}}, '{'{-25'd3664}}, '{'{25'd3331}}, '{'{-25'd466}}, '{'{25'd3398}}, '{'{25'd799}}, '{'{25'd733}}, '{'{-25'd5729}}, '{'{25'd1732}}, '{'{25'd1865}}, '{'{-25'd5929}}, '{'{25'd5463}}, '{'{-25'd5729}}, '{'{-25'd2065}}, '{'{25'd200}}, '{'{-25'd6862}}, '{'{25'd5263}}, '{'{25'd4130}}},
    '{'{'{-25'd4159}}, '{'{-25'd3866}}, '{'{25'd2109}}, '{'{25'd4452}}, '{'{25'd2577}}, '{'{-25'd3397}}, '{'{-25'd3514}}, '{'{-25'd7380}}, '{'{25'd4159}}, '{'{-25'd644}}, '{'{-25'd7380}}, '{'{25'd1406}}, '{'{-25'd2050}}, '{'{-25'd4569}}, '{'{25'd5975}}, '{'{25'd4217}}, '{'{25'd410}}, '{'{25'd4217}}, '{'{-25'd3866}}, '{'{25'd4217}}, '{'{-25'd4217}}, '{'{-25'd3339}}, '{'{-25'd4452}}, '{'{25'd351}}, '{'{-25'd5272}}, '{'{25'd3456}}, '{'{25'd3690}}, '{'{-25'd59}}, '{'{25'd3163}}, '{'{25'd4276}}, '{'{25'd2402}}, '{'{-25'd1640}}, '{'{25'd2519}}, '{'{-25'd2870}}, '{'{-25'd7087}}, '{'{-25'd3866}}, '{'{-25'd351}}, '{'{25'd1464}}, '{'{25'd879}}, '{'{25'd586}}, '{'{25'd3456}}, '{'{-25'd820}}, '{'{-25'd6677}}, '{'{-25'd5857}}, '{'{-25'd3983}}, '{'{25'd3104}}, '{'{-25'd4569}}, '{'{-25'd1816}}, '{'{25'd1581}}, '{'{-25'd2519}}, '{'{25'd117}}, '{'{25'd4510}}, '{'{25'd3924}}, '{'{25'd3632}}, '{'{25'd1640}}, '{'{-25'd4686}}, '{'{-25'd5330}}, '{'{25'd3983}}, '{'{-25'd1171}}, '{'{25'd3397}}, '{'{-25'd2167}}, '{'{-25'd2167}}, '{'{-25'd2694}}, '{'{-25'd4862}}},
    '{'{'{25'd4939}}, '{'{-25'd3669}}, '{'{25'd423}}, '{'{-25'd7197}}, '{'{-25'd1835}}, '{'{25'd3810}}, '{'{25'd1129}}, '{'{-25'd14677}}, '{'{-25'd3246}}, '{'{-25'd706}}, '{'{25'd2117}}, '{'{25'd2117}}, '{'{25'd565}}, '{'{-25'd8750}}, '{'{25'd6492}}, '{'{25'd1835}}, '{'{25'd3387}}, '{'{-25'd2823}}, '{'{25'd2823}}, '{'{-25'd4516}}, '{'{-25'd1976}}, '{'{25'd565}}, '{'{-25'd17641}}, '{'{-25'd10584}}, '{'{-25'd1270}}, '{'{-25'd282}}, '{'{25'd9032}}, '{'{-25'd4234}}, '{'{25'd2964}}, '{'{-25'd3387}}, '{'{-25'd2823}}, '{'{-25'd282}}, '{'{-25'd2964}}, '{'{25'd1694}}, '{'{-25'd1270}}, '{'{25'd3810}}, '{'{-25'd5927}}, '{'{-25'd1976}}, '{'{25'd2681}}, '{'{25'd2540}}, '{'{-25'd3528}}, '{'{-25'd4657}}, '{'{-25'd988}}, '{'{25'd17923}}, '{'{-25'd706}}, '{'{25'd3387}}, '{'{-25'd2823}}, '{'{-25'd5927}}, '{'{25'd3105}}, '{'{25'd8044}}, '{'{25'd7197}}, '{'{25'd0}}, '{'{25'd2258}}, '{'{25'd0}}, '{'{25'd8609}}, '{'{25'd423}}, '{'{25'd1129}}, '{'{-25'd3528}}, '{'{25'd1835}}, '{'{25'd3105}}, '{'{25'd3669}}, '{'{-25'd3669}}, '{'{-25'd2399}}, '{'{25'd3952}}},
    '{'{'{-25'd8089}}, '{'{25'd776}}, '{'{-25'd3878}}, '{'{-25'd7202}}, '{'{-25'd5872}}, '{'{25'd776}}, '{'{-25'd2216}}, '{'{25'd1551}}, '{'{-25'd4654}}, '{'{-25'd3435}}, '{'{25'd776}}, '{'{25'd2548}}, '{'{-25'd3878}}, '{'{25'd7978}}, '{'{-25'd111}}, '{'{25'd1108}}, '{'{25'd14072}}, '{'{-25'd3324}}, '{'{-25'd4764}}, '{'{25'd886}}, '{'{25'd3767}}, '{'{25'd5762}}, '{'{-25'd4100}}, '{'{25'd6205}}, '{'{-25'd886}}, '{'{25'd4764}}, '{'{25'd554}}, '{'{-25'd2548}}, '{'{-25'd4986}}, '{'{25'd3767}}, '{'{25'd5318}}, '{'{-25'd2216}}, '{'{25'd2327}}, '{'{-25'd4543}}, '{'{-25'd4432}}, '{'{25'd776}}, '{'{25'd1219}}, '{'{-25'd554}}, '{'{-25'd111}}, '{'{25'd5097}}, '{'{-25'd6205}}, '{'{25'd9086}}, '{'{-25'd1440}}, '{'{-25'd3767}}, '{'{-25'd776}}, '{'{25'd5872}}, '{'{-25'd3767}}, '{'{-25'd4100}}, '{'{-25'd2438}}, '{'{-25'd5208}}, '{'{-25'd3546}}, '{'{-25'd3102}}, '{'{-25'd6426}}, '{'{25'd5097}}, '{'{25'd3767}}, '{'{-25'd2770}}, '{'{25'd3324}}, '{'{25'd3102}}, '{'{25'd1551}}, '{'{-25'd4654}}, '{'{-25'd6981}}, '{'{-25'd7978}}, '{'{-25'd5540}}, '{'{25'd2881}}},
    '{'{'{-25'd1004}}, '{'{25'd91}}, '{'{-25'd2191}}, '{'{-25'd11231}}, '{'{25'd0}}, '{'{25'd730}}, '{'{-25'd2465}}, '{'{-25'd1187}}, '{'{25'd2557}}, '{'{25'd1278}}, '{'{25'd0}}, '{'{25'd2191}}, '{'{25'd1187}}, '{'{25'd3013}}, '{'{25'd730}}, '{'{-25'd3378}}, '{'{25'd11596}}, '{'{25'd3378}}, '{'{-25'd4292}}, '{'{25'd5205}}, '{'{-25'd3013}}, '{'{-25'd4931}}, '{'{25'd5113}}, '{'{-25'd5205}}, '{'{-25'd2557}}, '{'{-25'd5753}}, '{'{-25'd4565}}, '{'{25'd4657}}, '{'{25'd1004}}, '{'{25'd4018}}, '{'{-25'd2648}}, '{'{-25'd1278}}, '{'{25'd4018}}, '{'{-25'd5296}}, '{'{-25'd1552}}, '{'{-25'd3561}}, '{'{-25'd9222}}, '{'{25'd4931}}, '{'{-25'd1370}}, '{'{-25'd730}}, '{'{-25'd2557}}, '{'{25'd822}}, '{'{25'd4657}}, '{'{-25'd2831}}, '{'{25'd91}}, '{'{-25'd1644}}, '{'{25'd2374}}, '{'{25'd5022}}, '{'{-25'd5935}}, '{'{-25'd6574}}, '{'{-25'd3287}}, '{'{-25'd3105}}, '{'{25'd1644}}, '{'{-25'd5844}}, '{'{-25'd913}}, '{'{-25'd91}}, '{'{25'd3105}}, '{'{25'd1187}}, '{'{25'd9861}}, '{'{-25'd4292}}, '{'{25'd822}}, '{'{-25'd5296}}, '{'{-25'd1735}}, '{'{-25'd2009}}},
    '{'{'{-25'd4194}}, '{'{-25'd5266}}, '{'{-25'd585}}, '{'{25'd12386}}, '{'{25'd7119}}, '{'{-25'd1755}}, '{'{-25'd2438}}, '{'{25'd2341}}, '{'{25'd195}}, '{'{-25'd11020}}, '{'{-25'd4681}}, '{'{25'd975}}, '{'{-25'd1365}}, '{'{-25'd1073}}, '{'{25'd3511}}, '{'{-25'd1853}}, '{'{25'd9558}}, '{'{25'd1170}}, '{'{-25'd683}}, '{'{25'd3023}}, '{'{25'd4974}}, '{'{25'd1073}}, '{'{-25'd4779}}, '{'{25'd9362}}, '{'{-25'd2926}}, '{'{25'd3121}}, '{'{25'd2438}}, '{'{-25'd2146}}, '{'{-25'd293}}, '{'{-25'd3413}}, '{'{-25'd3218}}, '{'{-25'd2926}}, '{'{-25'd5559}}, '{'{-25'd878}}, '{'{25'd98}}, '{'{25'd1658}}, '{'{25'd8485}}, '{'{25'd4876}}, '{'{25'd585}}, '{'{-25'd10240}}, '{'{-25'd7705}}, '{'{-25'd1560}}, '{'{25'd3218}}, '{'{-25'd3316}}, '{'{25'd3706}}, '{'{-25'd1170}}, '{'{-25'd3901}}, '{'{-25'd3608}}, '{'{-25'd2438}}, '{'{-25'd1268}}, '{'{-25'd488}}, '{'{-25'd878}}, '{'{25'd3901}}, '{'{-25'd1365}}, '{'{25'd1268}}, '{'{-25'd1463}}, '{'{25'd5364}}, '{'{25'd7802}}, '{'{-25'd1853}}, '{'{25'd4389}}, '{'{-25'd3511}}, '{'{-25'd2438}}, '{'{-25'd5754}}, '{'{25'd5169}}},
    '{'{'{-25'd11847}}, '{'{-25'd4565}}, '{'{-25'd761}}, '{'{-25'd5978}}, '{'{25'd4239}}, '{'{-25'd3804}}, '{'{-25'd1848}}, '{'{25'd2608}}, '{'{-25'd3695}}, '{'{-25'd6086}}, '{'{-25'd3587}}, '{'{-25'd1739}}, '{'{25'd2608}}, '{'{-25'd3261}}, '{'{25'd217}}, '{'{25'd4673}}, '{'{-25'd5652}}, '{'{25'd435}}, '{'{-25'd1196}}, '{'{25'd6847}}, '{'{-25'd5217}}, '{'{-25'd3043}}, '{'{25'd5869}}, '{'{-25'd2391}}, '{'{25'd5108}}, '{'{-25'd1087}}, '{'{25'd3587}}, '{'{25'd978}}, '{'{-25'd2174}}, '{'{25'd1196}}, '{'{-25'd2391}}, '{'{-25'd3261}}, '{'{25'd6630}}, '{'{25'd5760}}, '{'{25'd326}}, '{'{-25'd11955}}, '{'{-25'd869}}, '{'{-25'd3369}}, '{'{25'd3152}}, '{'{-25'd109}}, '{'{25'd652}}, '{'{25'd5978}}, '{'{25'd2500}}, '{'{-25'd1522}}, '{'{25'd5869}}, '{'{25'd3913}}, '{'{-25'd543}}, '{'{25'd3478}}, '{'{25'd5434}}, '{'{25'd1087}}, '{'{-25'd5326}}, '{'{-25'd3804}}, '{'{25'd2174}}, '{'{-25'd2826}}, '{'{25'd3261}}, '{'{25'd2391}}, '{'{-25'd2174}}, '{'{25'd13803}}, '{'{-25'd1196}}, '{'{-25'd2391}}, '{'{-25'd2174}}, '{'{25'd2282}}, '{'{25'd1630}}, '{'{25'd761}}},
    '{'{'{-25'd863}}, '{'{-25'd2071}}, '{'{-25'd7078}}, '{'{-25'd9063}}, '{'{25'd3452}}, '{'{-25'd2417}}, '{'{25'd1640}}, '{'{25'd6991}}, '{'{-25'd1813}}, '{'{-25'd2071}}, '{'{-25'd5783}}, '{'{-25'd1899}}, '{'{25'd6732}}, '{'{25'd2330}}, '{'{-25'd3194}}, '{'{-25'd173}}, '{'{25'd5783}}, '{'{-25'd3452}}, '{'{25'd86}}, '{'{25'd3711}}, '{'{25'd2503}}, '{'{-25'd2589}}, '{'{-25'd2676}}, '{'{-25'd690}}, '{'{25'd3107}}, '{'{25'd2071}}, '{'{-25'd7164}}, '{'{25'd3711}}, '{'{25'd0}}, '{'{25'd6042}}, '{'{25'd2158}}, '{'{-25'd3280}}, '{'{25'd6560}}, '{'{-25'd3539}}, '{'{25'd3970}}, '{'{-25'd5092}}, '{'{25'd1122}}, '{'{25'd2503}}, '{'{-25'd1122}}, '{'{-25'd2417}}, '{'{-25'd10962}}, '{'{25'd6732}}, '{'{25'd5265}}, '{'{25'd259}}, '{'{-25'd3021}}, '{'{25'd0}}, '{'{-25'd2762}}, '{'{25'd1640}}, '{'{25'd86}}, '{'{-25'd6560}}, '{'{25'd949}}, '{'{25'd4661}}, '{'{-25'd2417}}, '{'{-25'd2330}}, '{'{-25'd949}}, '{'{25'd2330}}, '{'{-25'd3107}}, '{'{25'd6473}}, '{'{25'd8545}}, '{'{-25'd2158}}, '{'{25'd173}}, '{'{25'd3366}}, '{'{25'd5869}}, '{'{25'd2330}}},
    '{'{'{-25'd1389}}, '{'{-25'd2361}}, '{'{-25'd8888}}, '{'{25'd3750}}, '{'{-25'd278}}, '{'{25'd1111}}, '{'{25'd1389}}, '{'{25'd1389}}, '{'{-25'd4444}}, '{'{-25'd4444}}, '{'{-25'd5000}}, '{'{-25'd972}}, '{'{-25'd3194}}, '{'{25'd2916}}, '{'{25'd2500}}, '{'{-25'd3472}}, '{'{25'd17638}}, '{'{25'd4583}}, '{'{-25'd2361}}, '{'{25'd3750}}, '{'{25'd1944}}, '{'{-25'd1250}}, '{'{25'd1111}}, '{'{-25'd1250}}, '{'{25'd3889}}, '{'{-25'd3333}}, '{'{-25'd6111}}, '{'{-25'd2361}}, '{'{-25'd2916}}, '{'{25'd2222}}, '{'{-25'd3055}}, '{'{-25'd694}}, '{'{-25'd1389}}, '{'{25'd2778}}, '{'{25'd2916}}, '{'{-25'd6805}}, '{'{-25'd972}}, '{'{25'd3889}}, '{'{25'd1528}}, '{'{-25'd5555}}, '{'{-25'd14443}}, '{'{25'd3194}}, '{'{25'd4722}}, '{'{25'd7777}}, '{'{-25'd3472}}, '{'{25'd972}}, '{'{25'd3889}}, '{'{25'd1250}}, '{'{25'd2778}}, '{'{-25'd972}}, '{'{-25'd1250}}, '{'{-25'd2222}}, '{'{-25'd6527}}, '{'{-25'd2083}}, '{'{25'd4722}}, '{'{25'd972}}, '{'{-25'd2639}}, '{'{25'd9166}}, '{'{25'd3472}}, '{'{25'd3611}}, '{'{-25'd3055}}, '{'{25'd7638}}, '{'{25'd278}}, '{'{25'd556}}},
    '{'{'{25'd5749}}, '{'{-25'd7094}}, '{'{25'd5015}}, '{'{-25'd6361}}, '{'{-25'd5627}}, '{'{25'd2813}}, '{'{-25'd1101}}, '{'{25'd4648}}, '{'{25'd2324}}, '{'{-25'd5871}}, '{'{25'd2446}}, '{'{25'd3425}}, '{'{-25'd2079}}, '{'{25'd1835}}, '{'{-25'd3670}}, '{'{25'd5871}}, '{'{25'd10642}}, '{'{-25'd1468}}, '{'{25'd3180}}, '{'{-25'd4281}}, '{'{-25'd4648}}, '{'{25'd1712}}, '{'{-25'd2446}}, '{'{-25'd2446}}, '{'{-25'd1835}}, '{'{-25'd367}}, '{'{25'd4281}}, '{'{25'd1346}}, '{'{-25'd4037}}, '{'{25'd1101}}, '{'{25'd5504}}, '{'{25'd979}}, '{'{25'd3670}}, '{'{-25'd2936}}, '{'{-25'd1468}}, '{'{-25'd5749}}, '{'{25'd9052}}, '{'{-25'd3058}}, '{'{25'd979}}, '{'{-25'd6238}}, '{'{25'd3425}}, '{'{25'd15534}}, '{'{25'd1346}}, '{'{-25'd2813}}, '{'{25'd489}}, '{'{25'd1468}}, '{'{25'd3180}}, '{'{25'd2569}}, '{'{-25'd1101}}, '{'{25'd734}}, '{'{25'd0}}, '{'{25'd856}}, '{'{-25'd7951}}, '{'{-25'd3547}}, '{'{25'd5749}}, '{'{-25'd3670}}, '{'{25'd2446}}, '{'{25'd2691}}, '{'{-25'd8073}}, '{'{-25'd2446}}, '{'{-25'd5015}}, '{'{-25'd10764}}, '{'{25'd122}}, '{'{-25'd3425}}},
    '{'{'{25'd2021}}, '{'{-25'd1235}}, '{'{25'd2358}}, '{'{-25'd4492}}, '{'{25'd561}}, '{'{25'd4829}}, '{'{25'd1011}}, '{'{25'd4155}}, '{'{-25'd2695}}, '{'{-25'd5839}}, '{'{-25'd6064}}, '{'{-25'd3594}}, '{'{25'd225}}, '{'{25'd5053}}, '{'{25'd4043}}, '{'{25'd6289}}, '{'{25'd14262}}, '{'{25'd2920}}, '{'{-25'd5053}}, '{'{25'd561}}, '{'{-25'd4380}}, '{'{25'd2358}}, '{'{25'd3257}}, '{'{-25'd7299}}, '{'{25'd3481}}, '{'{-25'd4716}}, '{'{-25'd5053}}, '{'{25'd3032}}, '{'{-25'd3594}}, '{'{-25'd337}}, '{'{25'd2471}}, '{'{25'd2583}}, '{'{25'd5727}}, '{'{-25'd2471}}, '{'{25'd112}}, '{'{25'd674}}, '{'{25'd3369}}, '{'{-25'd5053}}, '{'{-25'd5615}}, '{'{-25'd5390}}, '{'{-25'd1011}}, '{'{25'd898}}, '{'{-25'd1684}}, '{'{25'd0}}, '{'{-25'd3481}}, '{'{25'd1235}}, '{'{25'd3706}}, '{'{25'd5278}}, '{'{25'd4492}}, '{'{25'd1011}}, '{'{25'd6401}}, '{'{25'd1123}}, '{'{-25'd3818}}, '{'{-25'd1123}}, '{'{25'd337}}, '{'{-25'd4492}}, '{'{-25'd2246}}, '{'{25'd3369}}, '{'{25'd2358}}, '{'{-25'd6626}}, '{'{-25'd5166}}, '{'{25'd2807}}, '{'{25'd4829}}, '{'{-25'd1909}}},
    '{'{'{25'd3141}}, '{'{-25'd6374}}, '{'{-25'd4342}}, '{'{25'd6744}}, '{'{25'd7945}}, '{'{25'd1016}}, '{'{25'd1848}}, '{'{-25'd2217}}, '{'{25'd3603}}, '{'{-25'd3141}}, '{'{-25'd2494}}, '{'{25'd4342}}, '{'{-25'd370}}, '{'{-25'd2402}}, '{'{25'd6559}}, '{'{25'd1293}}, '{'{25'd9146}}, '{'{25'd1848}}, '{'{25'd3326}}, '{'{-25'd3603}}, '{'{25'd1663}}, '{'{-25'd3788}}, '{'{-25'd6005}}, '{'{25'd554}}, '{'{25'd4157}}, '{'{-25'd2032}}, '{'{25'd1848}}, '{'{-25'd4804}}, '{'{-25'd647}}, '{'{-25'd3233}}, '{'{-25'd2956}}, '{'{-25'd4804}}, '{'{-25'd4619}}, '{'{25'd3880}}, '{'{-25'd4342}}, '{'{-25'd2402}}, '{'{25'd2309}}, '{'{25'd2587}}, '{'{-25'd554}}, '{'{-25'd277}}, '{'{-25'd11178}}, '{'{25'd11732}}, '{'{-25'd3233}}, '{'{25'd4342}}, '{'{25'd2402}}, '{'{25'd4434}}, '{'{25'd1478}}, '{'{-25'd5081}}, '{'{25'd0}}, '{'{-25'd8776}}, '{'{25'd4619}}, '{'{-25'd2125}}, '{'{25'd0}}, '{'{25'd4988}}, '{'{25'd1478}}, '{'{-25'd2679}}, '{'{-25'd3049}}, '{'{25'd3049}}, '{'{-25'd2771}}, '{'{-25'd185}}, '{'{-25'd9330}}, '{'{25'd3233}}, '{'{25'd3418}}, '{'{-25'd2587}}},
    '{'{'{-25'd10274}}, '{'{-25'd5618}}, '{'{-25'd1364}}, '{'{-25'd6341}}, '{'{25'd1284}}, '{'{-25'd3853}}, '{'{-25'd4414}}, '{'{25'd4414}}, '{'{-25'd2488}}, '{'{-25'd4976}}, '{'{25'd883}}, '{'{-25'd963}}, '{'{25'd5538}}, '{'{25'd0}}, '{'{-25'd1605}}, '{'{-25'd2649}}, '{'{25'd4896}}, '{'{-25'd3130}}, '{'{25'd2809}}, '{'{-25'd1445}}, '{'{-25'd3130}}, '{'{-25'd2729}}, '{'{25'd3853}}, '{'{-25'd4495}}, '{'{25'd4254}}, '{'{-25'd3933}}, '{'{25'd3130}}, '{'{25'd3532}}, '{'{25'd3853}}, '{'{-25'd2247}}, '{'{25'd1766}}, '{'{-25'd2167}}, '{'{-25'd3692}}, '{'{-25'd1204}}, '{'{25'd1204}}, '{'{-25'd1605}}, '{'{-25'd80}}, '{'{25'd2488}}, '{'{25'd2328}}, '{'{-25'd7545}}, '{'{-25'd3933}}, '{'{25'd10193}}, '{'{25'd4254}}, '{'{25'd2809}}, '{'{25'd2649}}, '{'{25'd4334}}, '{'{25'd5217}}, '{'{-25'd80}}, '{'{-25'd4896}}, '{'{-25'd4896}}, '{'{25'd4334}}, '{'{25'd4013}}, '{'{-25'd8347}}, '{'{-25'd4174}}, '{'{25'd1124}}, '{'{-25'd2889}}, '{'{25'd6100}}, '{'{25'd6501}}, '{'{25'd10193}}, '{'{25'd321}}, '{'{25'd0}}, '{'{-25'd7464}}, '{'{25'd2809}}, '{'{-25'd1204}}},
    '{'{'{-25'd4062}}, '{'{-25'd5109}}, '{'{-25'd6216}}, '{'{25'd2216}}, '{'{-25'd2400}}, '{'{25'd3754}}, '{'{25'd5786}}, '{'{-25'd3878}}, '{'{-25'd800}}, '{'{-25'd800}}, '{'{-25'd2585}}, '{'{25'd4555}}, '{'{25'd3139}}, '{'{25'd308}}, '{'{25'd3570}}, '{'{-25'd1600}}, '{'{-25'd185}}, '{'{-25'd4431}}, '{'{-25'd2770}}, '{'{25'd4862}}, '{'{25'd5047}}, '{'{25'd800}}, '{'{25'd4678}}, '{'{-25'd7878}}, '{'{-25'd2647}}, '{'{25'd1662}}, '{'{-25'd1354}}, '{'{-25'd1046}}, '{'{-25'd2277}}, '{'{25'd5355}}, '{'{25'd123}}, '{'{25'd3693}}, '{'{-25'd5170}}, '{'{25'd308}}, '{'{-25'd1416}}, '{'{25'd2831}}, '{'{25'd1970}}, '{'{-25'd1662}}, '{'{-25'd4185}}, '{'{-25'd6340}}, '{'{-25'd1908}}, '{'{25'd2585}}, '{'{-25'd3754}}, '{'{25'd2647}}, '{'{25'd800}}, '{'{25'd1046}}, '{'{-25'd1723}}, '{'{-25'd2339}}, '{'{25'd2831}}, '{'{-25'd5478}}, '{'{25'd3385}}, '{'{25'd5416}}, '{'{25'd1662}}, '{'{-25'd2647}}, '{'{25'd2523}}, '{'{-25'd3016}}, '{'{-25'd1723}}, '{'{25'd6340}}, '{'{25'd4801}}, '{'{-25'd985}}, '{'{-25'd4924}}, '{'{-25'd308}}, '{'{-25'd862}}, '{'{-25'd3139}}},
    '{'{'{-25'd2070}}, '{'{25'd966}}, '{'{25'd2760}}, '{'{25'd8350}}, '{'{25'd966}}, '{'{25'd5107}}, '{'{25'd5797}}, '{'{25'd2553}}, '{'{-25'd3312}}, '{'{-25'd6073}}, '{'{25'd897}}, '{'{25'd1242}}, '{'{-25'd69}}, '{'{-25'd3105}}, '{'{-25'd1104}}, '{'{-25'd3933}}, '{'{25'd8764}}, '{'{-25'd828}}, '{'{25'd1035}}, '{'{-25'd414}}, '{'{-25'd3105}}, '{'{-25'd2139}}, '{'{-25'd1449}}, '{'{-25'd4486}}, '{'{-25'd5314}}, '{'{-25'd1380}}, '{'{-25'd897}}, '{'{25'd0}}, '{'{25'd621}}, '{'{-25'd3588}}, '{'{-25'd3795}}, '{'{25'd1518}}, '{'{25'd1242}}, '{'{25'd759}}, '{'{-25'd2415}}, '{'{-25'd4071}}, '{'{25'd5314}}, '{'{25'd2622}}, '{'{-25'd2829}}, '{'{-25'd7039}}, '{'{-25'd5935}}, '{'{-25'd2277}}, '{'{25'd3381}}, '{'{25'd2553}}, '{'{25'd5245}}, '{'{-25'd345}}, '{'{25'd2139}}, '{'{25'd7315}}, '{'{25'd6349}}, '{'{-25'd3795}}, '{'{25'd1380}}, '{'{25'd4209}}, '{'{-25'd3864}}, '{'{-25'd4900}}, '{'{-25'd552}}, '{'{25'd2001}}, '{'{-25'd207}}, '{'{25'd4693}}, '{'{25'd552}}, '{'{-25'd3657}}, '{'{25'd3105}}, '{'{25'd4831}}, '{'{-25'd2967}}, '{'{-25'd2070}}},
    '{'{'{25'd5358}}, '{'{-25'd3006}}, '{'{-25'd1699}}, '{'{-25'd2091}}, '{'{-25'd4574}}, '{'{25'd4574}}, '{'{25'd523}}, '{'{25'd6926}}, '{'{-25'd3006}}, '{'{-25'd1960}}, '{'{25'd2614}}, '{'{-25'd2352}}, '{'{25'd5358}}, '{'{-25'd3267}}, '{'{-25'd6926}}, '{'{25'd6403}}, '{'{25'd16597}}, '{'{-25'd915}}, '{'{-25'd2352}}, '{'{25'd1830}}, '{'{-25'd1438}}, '{'{-25'd653}}, '{'{-25'd523}}, '{'{-25'd6011}}, '{'{-25'd4835}}, '{'{25'd3659}}, '{'{25'd4835}}, '{'{25'd3659}}, '{'{25'd1830}}, '{'{-25'd1307}}, '{'{25'd7057}}, '{'{-25'd5097}}, '{'{25'd2614}}, '{'{25'd3921}}, '{'{25'd1568}}, '{'{-25'd4835}}, '{'{25'd7580}}, '{'{-25'd1176}}, '{'{-25'd3921}}, '{'{25'd915}}, '{'{-25'd10455}}, '{'{25'd4835}}, '{'{-25'd4966}}, '{'{25'd3267}}, '{'{-25'd3267}}, '{'{-25'd4051}}, '{'{25'd6011}}, '{'{-25'd1699}}, '{'{-25'd7188}}, '{'{25'd3790}}, '{'{-25'd3790}}, '{'{25'd1045}}, '{'{-25'd9540}}, '{'{25'd915}}, '{'{-25'd2091}}, '{'{25'd1307}}, '{'{25'd2222}}, '{'{25'd11762}}, '{'{-25'd10063}}, '{'{25'd4182}}, '{'{-25'd4835}}, '{'{25'd1045}}, '{'{-25'd1307}}, '{'{25'd5227}}}
};
