localparam bit signed [0:146][7:0] Input1 = '{-86, 59, 95, -74, 73, -13, 51, -46, -105, -45, -103, -71, 69, -39, -83, -17, -40, 51, -69, 44, 26, -8, -11, 43, -7, 32, -98, 14, -57, -32, 61, -127, 118, 47, -4, -19, -10, 43, 90, -113, -60, 74, -43, 39, -22, 107, -34, 86, -128, -47, 58, -116, 91, -85, 54, -3, 47, -106, -97, -12, -94, 98, -86, -60, -6, -66, -92, -45, 44, 81, 112, -17, 70, -122, 48, 9, -100, -51, 56, 9, 85, -62, -119, -18, 120, 36, -100, 116, -64, 74, -4, 13, 107, -126, 37, 71, -41, 94, 81, -125, -17, 98, -48, 115, -46, -78, 61, 106, 82, -100, -93, -75, -102, -15, -25, -86, -82, 69, -100, -1, 43, -45, -66, -54, 74, 9, 91, 99, -53, -32, 38, -97, 115, 22, -2, -37, -71, -107, 97, -67, 108, -87, -13, -21, -29, 41, 122};
