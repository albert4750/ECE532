logic signed [15:0] layer3_weight[3][8][3][3] = '{
    '{
        '{'{9435, 21122, -27768}, '{21576, -2343, 6438}, '{-31180, -287, 18776}},
        '{'{15679, -21611, 31236}, '{18847, -23821, 14539}, '{-1371, -2297, -12650}},
        '{'{28284, -6870, 22715}, '{-21793, 16694, -10295}, '{-16525, -19021, -5550}},
        '{'{-4329, -17325, -10471}, '{-10439, 23749, 22873}, '{16685, 15727, -2472}},
        '{'{-6221, -31429, -14420}, '{-15206, 3704, 19061}, '{31659, 21113, -7776}},
        '{'{-6370, -26994, -12985}, '{28768, -14659, 513}, '{3574, -18001, -25220}},
        '{'{18797, 11382, -9045}, '{-13862, 25615, 8004}, '{-15158, -10155, -4441}},
        '{'{106, -25109, 13918}, '{32214, -28416, 9809}, '{19642, -5108, 21723}}
    },
    '{
        '{'{-17621, -27722, -1667}, '{-7761, -23786, 15135}, '{-20108, 15394, 26594}},
        '{'{28458, -29372, 3962}, '{17214, 3876, -4269}, '{-5972, -23855, -22288}},
        '{'{-17041, 8390, -7930}, '{-29264, 30089, 24092}, '{20557, 30392, -30327}},
        '{'{469, 26434, 14857}, '{29806, 7160, -31580}, '{8476, 22004, -17344}},
        '{'{-15414, 13180, -2931}, '{-789, 26114, -30299}, '{-9273, 7255, 1758}},
        '{'{4049, 26115, -16273}, '{-18462, -25776, -30989}, '{-28078, -11470, 18365}},
        '{'{-30230, 29650, -20452}, '{1827, 24885, 12058}, '{-29327, -27289, -27094}},
        '{'{28462, -3899, 23068}, '{-8065, 24747, -23469}, '{20542, -1206, 11466}}
    },
    '{
        '{'{23177, -15141, -27933}, '{15179, -13472, 28838}, '{22559, -20749, -8298}},
        '{'{-29314, -2213, 5945}, '{23573, 28385, -28867}, '{-532, 3881, -1677}},
        '{'{-11413, 26979, 31913}, '{-5894, -24937, -8963}, '{-29976, 5940, -32489}},
        '{'{-23430, 20296, -20951}, '{19693, -19652, -31953}, '{9871, 29732, -26687}},
        '{'{2654, -22555, -15574}, '{-8450, 512, -45}, '{19334, -27939, 3139}},
        '{'{-28385, -29923, -26608}, '{-6205, -1766, -12291}, '{25862, -12055, 11749}},
        '{'{-12021, -29359, -21705}, '{4989, -23253, 6467}, '{-19948, 12763, -32257}},
        '{'{19063, 13788, -28402}, '{-16114, -6064, 15843}, '{-32321, 4469, 16102}}
    }
};
