localparam bit signed [0:146][7:0] Input3 = '{-44, -107, -9, -101, 26, 89, 64, -18, 3, -75, -91, -121, -8, -48, 75, 11, 108, 2, -74, -123, -111, 122, -3, -50, 5, -50, -47, 105, -18, -20, -98, -30, -125, 0, -35, -84, 44, 108, -1, -13, 61, 126, -128, -111, 29, -37, 34, 114, 115, 100, 59, -107, -65, 94, 120, -27, 17, -90, 79, 1, 15, 105, 86, 109, -111, 108, 53, 22, 77, -14, 47, 66, -117, 9, 114, -88, 54, 51, -81, -124, 10, 113, 126, 6, -10, 44, -56, 8, 72, 108, 101, -110, -126, 69, 93, 121, 101, -28, -22, 29, 27, 17, 58, 11, -79, -56, -40, -125, -16, -117, -71, 50, 15, 57, 3, -10, 100, 60, 39, 126, 85, 29, 53, -61, -72, 75, -9, -49, -83, -38, -49, 97, -117, 119, 5, 30, 58, -60, -69, -96, -91, 43, -3, -68, -83, -99, 122};
