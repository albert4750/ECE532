logic signed [7:0] convolve6_weight[4][8][3][3] = '{
    '{
        '{'{112, 66, 47}, '{-111, -108, 38}, '{-64, 6, 108}},
        '{'{22, -49, -54}, '{34, 40, 38}, '{118, 21, -94}},
        '{'{-11, 32, 42}, '{-1, -84, -29}, '{-87, 121, -25}},
        '{'{27, 123, -80}, '{-1, 10, -60}, '{-111, -125, -27}},
        '{'{-34, 87, -99}, '{-26, -5, 30}, '{75, 66, 93}},
        '{'{-68, 7, 51}, '{116, -55, 87}, '{64, 112, 17}},
        '{'{40, 115, -107}, '{-34, 26, 15}, '{112, -111, -118}},
        '{'{17, 3, 103}, '{-55, -99, 67}, '{71, 80, 98}}
    },
    '{
        '{'{4, 61, -38}, '{-28, 6, -96}, '{-47, -9, -10}},
        '{'{117, -91, -9}, '{-101, -77, -50}, '{59, -42, -33}},
        '{'{-120, -72, -99}, '{28, 95, 34}, '{58, -1, -2}},
        '{'{81, 92, -17}, '{16, 72, -69}, '{119, 108, -121}},
        '{'{12, -96, 84}, '{107, -53, 93}, '{-88, -128, 84}},
        '{'{-19, -36, 77}, '{37, 47, -67}, '{-25, 50, -60}},
        '{'{110, 76, 57}, '{-9, 101, 112}, '{4, -23, -92}},
        '{'{-48, 82, 37}, '{94, -11, 110}, '{-93, 48, 0}}
    },
    '{
        '{'{-79, 57, -119}, '{-78, 97, 48}, '{113, -116, 70}},
        '{'{-4, 115, 36}, '{-29, -26, -92}, '{-98, -14, 19}},
        '{'{38, 44, -93}, '{-114, -99, 51}, '{-68, 120, -47}},
        '{'{-61, -99, 27}, '{3, -95, 117}, '{51, -10, 27}},
        '{'{100, -72, -107}, '{39, 106, -54}, '{-99, 113, 29}},
        '{'{61, -70, -104}, '{-14, -112, 64}, '{-28, 98, -5}},
        '{'{-115, -127, 123}, '{-126, -62, 19}, '{116, 122, 76}},
        '{'{30, -89, 85}, '{-51, 49, -102}, '{-13, 12, 113}}
    },
    '{
        '{'{64, -127, 36}, '{-118, -22, -96}, '{126, -100, 58}},
        '{'{66, 92, -63}, '{77, -45, -81}, '{-47, 36, 71}},
        '{'{-75, 70, 9}, '{-113, -110, 29}, '{53, 60, -86}},
        '{'{82, 2, -99}, '{17, -93, -8}, '{-109, 16, -105}},
        '{'{12, -29, -19}, '{56, 66, -108}, '{3, -47, 44}},
        '{'{-90, -86, 74}, '{-91, -22, -88}, '{-17, -101, 4}},
        '{'{51, 22, 37}, '{-93, -98, -121}, '{88, -40, 111}},
        '{'{15, 10, 19}, '{-51, 103, -72}, '{101, 103, 18}}
    }
};
