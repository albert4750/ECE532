localparam bit signed [0:7][36:0] Bias1 = '{37'd0, 37'd0, 37'd0, 37'd0, 37'd0, 37'd0, 37'd0, 37'd0};
