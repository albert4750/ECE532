localparam bit signed [0:31][0:63][0:0][0:0][24:0] Weight2 = '{
    '{'{'{-25'd1576991}}, '{'{25'd1506902}}, '{'{-25'd946195}}, '{'{-25'd665841}}, '{'{-25'd946195}}, '{'{25'd350442}}, '{'{25'd420531}}, '{'{25'd0}}, '{'{25'd315398}}, '{'{-25'd490619}}, '{'{-25'd1366725}}, '{'{25'd245310}}, '{'{25'd1787256}}, '{'{25'd735929}}, '{'{-25'd700885}}, '{'{25'd700885}}, '{'{25'd1296637}}, '{'{25'd1051327}}, '{'{25'd1156460}}, '{'{25'd175221}}, '{'{-25'd4485663}}, '{'{-25'd630796}}, '{'{25'd1016283}}, '{'{-25'd420531}}, '{'{25'd1366725}}, '{'{-25'd560708}}, '{'{-25'd560708}}, '{'{-25'd1541947}}, '{'{-25'd525664}}, '{'{-25'd700885}}, '{'{-25'd245310}}, '{'{25'd1086372}}, '{'{25'd70088}}, '{'{25'd280354}}, '{'{25'd560708}}, '{'{-25'd1261593}}, '{'{-25'd1752212}}, '{'{-25'd630796}}, '{'{-25'd1752212}}, '{'{25'd490619}}, '{'{-25'd911150}}, '{'{-25'd175221}}, '{'{25'd35044}}, '{'{25'd946195}}, '{'{25'd1296637}}, '{'{-25'd70088}}, '{'{25'd1471858}}, '{'{-25'd700885}}, '{'{-25'd946195}}, '{'{25'd1612035}}, '{'{-25'd35044}}, '{'{25'd981239}}, '{'{25'd981239}}, '{'{25'd210265}}, '{'{-25'd455575}}, '{'{-25'd1541947}}, '{'{25'd770973}}, '{'{25'd1436814}}, '{'{25'd280354}}, '{'{-25'd1051327}}, '{'{-25'd981239}}, '{'{25'd420531}}, '{'{25'd1261593}}, '{'{25'd1331681}}},
    '{'{'{25'd190454}}, '{'{-25'd269810}}, '{'{25'd730074}}, '{'{25'd1618859}}, '{'{-25'd396779}}, '{'{-25'd1031626}}, '{'{-25'd1650601}}, '{'{-25'd618975}}, '{'{25'd1380791}}, '{'{-25'd603104}}, '{'{-25'd190454}}, '{'{-25'd1507761}}, '{'{25'd301552}}, '{'{25'd317423}}, '{'{25'd412650}}, '{'{-25'd888785}}, '{'{-25'd365037}}, '{'{25'd745945}}, '{'{25'd1333178}}, '{'{25'd650718}}, '{'{25'd825301}}, '{'{25'd333294}}, '{'{-25'd571362}}, '{'{25'd603104}}, '{'{25'd47613}}, '{'{25'd285681}}, '{'{25'd1253822}}, '{'{-25'd1587116}}, '{'{-25'd698331}}, '{'{-25'd1158595}}, '{'{-25'd285681}}, '{'{25'd682460}}, '{'{25'd539620}}, '{'{25'd1650601}}, '{'{25'd825301}}, '{'{25'd1174466}}, '{'{-25'd301552}}, '{'{25'd1079239}}, '{'{-25'd634847}}, '{'{-25'd1174466}}, '{'{-25'd1190337}}, '{'{25'd1412534}}, '{'{-25'd380908}}, '{'{25'd777687}}, '{'{25'd1523632}}, '{'{25'd365037}}, '{'{25'd1206208}}, '{'{-25'd285681}}, '{'{-25'd1015754}}, '{'{25'd349166}}, '{'{25'd666589}}, '{'{25'd1761699}}, '{'{25'd793558}}, '{'{-25'd460264}}, '{'{-25'd2031509}}, '{'{-25'd1587116}}, '{'{25'd603104}}, '{'{25'd1793442}}, '{'{-25'd15871}}, '{'{-25'd174583}}, '{'{-25'd1539503}}, '{'{-25'd1110981}}, '{'{25'd95227}}, '{'{-25'd317423}}},
    '{'{'{25'd232888}}, '{'{25'd873331}}, '{'{-25'd1106219}}, '{'{25'd1164441}}, '{'{25'd1863105}}, '{'{25'd1571995}}, '{'{-25'd1921327}}, '{'{25'd640442}}, '{'{25'd1630217}}, '{'{-25'd1688439}}, '{'{25'd0}}, '{'{25'd465776}}, '{'{25'd0}}, '{'{-25'd7452421}}, '{'{-25'd640442}}, '{'{25'd815109}}, '{'{-25'd1047997}}, '{'{-25'd1571995}}, '{'{-25'd698664}}, '{'{-25'd2911102}}, '{'{25'd1455551}}, '{'{-25'd2154215}}, '{'{25'd174666}}, '{'{-25'd1164441}}, '{'{25'd1047997}}, '{'{25'd1746661}}, '{'{-25'd1746661}}, '{'{25'd349332}}, '{'{25'd1164441}}, '{'{25'd3726210}}, '{'{25'd1339107}}, '{'{25'd815109}}, '{'{25'd698664}}, '{'{-25'd1047997}}, '{'{-25'd989775}}, '{'{25'd1164441}}, '{'{25'd465776}}, '{'{25'd698664}}, '{'{-25'd2037771}}, '{'{-25'd407554}}, '{'{-25'd1339107}}, '{'{25'd407554}}, '{'{25'd1222663}}, '{'{25'd1280885}}, '{'{25'd232888}}, '{'{-25'd1513773}}, '{'{-25'd1455551}}, '{'{-25'd1047997}}, '{'{25'd407554}}, '{'{25'd582220}}, '{'{25'd232888}}, '{'{-25'd465776}}, '{'{25'd349332}}, '{'{25'd465776}}, '{'{25'd1047997}}, '{'{-25'd1280885}}, '{'{-25'd815109}}, '{'{-25'd1397329}}, '{'{-25'd116444}}, '{'{25'd116444}}, '{'{25'd640442}}, '{'{-25'd1106219}}, '{'{-25'd1397329}}, '{'{25'd349332}}},
    '{'{'{-25'd28634}}, '{'{25'd773109}}, '{'{25'd372238}}, '{'{-25'd214752}}, '{'{-25'd816059}}, '{'{-25'd744475}}, '{'{-25'd486772}}, '{'{25'd1102396}}, '{'{-25'd973545}}, '{'{25'd1446000}}, '{'{25'd1589168}}, '{'{-25'd42950}}, '{'{-25'd601307}}, '{'{25'd1102396}}, '{'{-25'd744475}}, '{'{-25'd1546218}}, '{'{-25'd1360099}}, '{'{25'd744475}}, '{'{-25'd157485}}, '{'{25'd343604}}, '{'{25'd1460317}}, '{'{-25'd1331465}}, '{'{-25'd186119}}, '{'{25'd200436}}, '{'{-25'd1302832}}, '{'{25'd1016495}}, '{'{-25'd787426}}, '{'{25'd1188297}}, '{'{-25'd959228}}, '{'{-25'd1732337}}, '{'{-25'd1517584}}, '{'{25'd429505}}, '{'{25'd1818238}}, '{'{25'd601307}}, '{'{-25'd773109}}, '{'{25'd157485}}, '{'{-25'd1431683}}, '{'{25'd1560535}}, '{'{25'd544040}}, '{'{25'd501089}}, '{'{25'd1030812}}, '{'{25'd1789604}}, '{'{25'd1732337}}, '{'{-25'd458139}}, '{'{-25'd429505}}, '{'{25'd243386}}, '{'{-25'd300653}}, '{'{25'd1703703}}, '{'{25'd1374416}}, '{'{25'd730158}}, '{'{-25'd1603485}}, '{'{-25'd415188}}, '{'{-25'd515406}}, '{'{25'd1431683}}, '{'{25'd42950}}, '{'{-25'd243386}}, '{'{25'd773109}}, '{'{25'd443822}}, '{'{25'd1617802}}, '{'{-25'd544040}}, '{'{25'd42950}}, '{'{25'd1216931}}, '{'{-25'd1460317}}, '{'{25'd787426}}},
    '{'{'{25'd388619}}, '{'{25'd340042}}, '{'{-25'd906778}}, '{'{25'd2056444}}, '{'{25'd1133473}}, '{'{25'd939163}}, '{'{25'd906778}}, '{'{25'd1230628}}, '{'{-25'd744854}}, '{'{-25'd323849}}, '{'{-25'd1457322}}, '{'{-25'd955356}}, '{'{25'd2056444}}, '{'{-25'd242887}}, '{'{-25'd1182050}}, '{'{-25'd890586}}, '{'{25'd32385}}, '{'{25'd485774}}, '{'{25'd32385}}, '{'{-25'd1279205}}, '{'{-25'd242887}}, '{'{25'd1554477}}, '{'{25'd97155}}, '{'{25'd680084}}, '{'{-25'd1441130}}, '{'{-25'd874393}}, '{'{-25'd1473515}}, '{'{25'd1101088}}, '{'{-25'd1554477}}, '{'{25'd1052511}}, '{'{25'd1959289}}, '{'{-25'd80962}}, '{'{-25'd1441130}}, '{'{-25'd340042}}, '{'{-25'd858201}}, '{'{25'd1052511}}, '{'{25'd615314}}, '{'{-25'd1182050}}, '{'{25'd1975481}}, '{'{-25'd16192}}, '{'{25'd1101088}}, '{'{-25'd1182050}}, '{'{25'd793431}}, '{'{-25'd955356}}, '{'{25'd404812}}, '{'{25'd663891}}, '{'{25'd323849}}, '{'{25'd1311590}}, '{'{-25'd647699}}, '{'{-25'd356234}}, '{'{25'd1214435}}, '{'{-25'd80962}}, '{'{25'd1376360}}, '{'{25'd615314}}, '{'{25'd939163}}, '{'{25'd178117}}, '{'{25'd469582}}, '{'{-25'd1635439}}, '{'{25'd1522092}}, '{'{-25'd340042}}, '{'{25'd80962}}, '{'{25'd1716402}}, '{'{25'd437197}}, '{'{25'd1230628}}},
    '{'{'{25'd94806}}, '{'{-25'd94806}}, '{'{-25'd995467}}, '{'{25'd1896128}}, '{'{25'd616242}}, '{'{-25'd1611709}}, '{'{25'd1327290}}, '{'{-25'd1516903}}, '{'{-25'd521435}}, '{'{-25'd1469499}}, '{'{-25'd900661}}, '{'{-25'd331822}}, '{'{25'd6020207}}, '{'{25'd2133144}}, '{'{25'd1422096}}, '{'{25'd379226}}, '{'{-25'd568838}}, '{'{-25'd47403}}, '{'{-25'd189613}}, '{'{-25'd189613}}, '{'{-25'd3887063}}, '{'{25'd711048}}, '{'{25'd4835127}}, '{'{25'd1327290}}, '{'{-25'd2701983}}, '{'{25'd1090274}}, '{'{25'd1848725}}, '{'{-25'd284419}}, '{'{-25'd616242}}, '{'{-25'd711048}}, '{'{-25'd474032}}, '{'{-25'd711048}}, '{'{25'd3223418}}, '{'{-25'd237016}}, '{'{-25'd1753919}}, '{'{-25'd1801322}}, '{'{25'd142210}}, '{'{-25'd1753919}}, '{'{25'd1327290}}, '{'{25'd568838}}, '{'{25'd284419}}, '{'{25'd1706515}}, '{'{25'd1279887}}, '{'{25'd1469499}}, '{'{25'd1327290}}, '{'{-25'd853258}}, '{'{25'd47403}}, '{'{-25'd900661}}, '{'{25'd331822}}, '{'{25'd948064}}, '{'{25'd1232483}}, '{'{25'd2180548}}, '{'{-25'd1137677}}, '{'{-25'd1327290}}, '{'{-25'd1374693}}, '{'{-25'd948064}}, '{'{-25'd1042871}}, '{'{25'd0}}, '{'{25'd1943532}}, '{'{25'd663645}}, '{'{-25'd142210}}, '{'{25'd142210}}, '{'{25'd1327290}}, '{'{-25'd426629}}},
    '{'{'{-25'd858760}}, '{'{-25'd143127}}, '{'{25'd477089}}, '{'{-25'd572507}}, '{'{-25'd858760}}, '{'{-25'd1669811}}, '{'{-25'd858760}}, '{'{25'd1240431}}, '{'{25'd667924}}, '{'{-25'd1001887}}, '{'{-25'd1192722}}, '{'{-25'd1478975}}, '{'{25'd620215}}, '{'{25'd1240431}}, '{'{-25'd1622102}}, '{'{25'd1097304}}, '{'{-25'd286253}}, '{'{25'd1192722}}, '{'{-25'd620215}}, '{'{-25'd954178}}, '{'{-25'd1717520}}, '{'{25'd2337735}}, '{'{-25'd381671}}, '{'{25'd238544}}, '{'{25'd190836}}, '{'{-25'd1192722}}, '{'{-25'd1478975}}, '{'{-25'd286253}}, '{'{25'd0}}, '{'{25'd6059028}}, '{'{-25'd1526684}}, '{'{-25'd1956064}}, '{'{25'd1431267}}, '{'{25'd954178}}, '{'{25'd1145013}}, '{'{-25'd95418}}, '{'{-25'd381671}}, '{'{-25'd1097304}}, '{'{25'd2528571}}, '{'{-25'd1335849}}, '{'{25'd4866306}}, '{'{25'd190836}}, '{'{25'd1860646}}, '{'{25'd1335849}}, '{'{-25'd1622102}}, '{'{-25'd1383558}}, '{'{-25'd1049595}}, '{'{-25'd333962}}, '{'{25'd190836}}, '{'{25'd1240431}}, '{'{25'd2433153}}, '{'{25'd1860646}}, '{'{25'd1097304}}, '{'{-25'd715633}}, '{'{25'd47709}}, '{'{25'd1049595}}, '{'{-25'd811051}}, '{'{-25'd1288140}}, '{'{-25'd667924}}, '{'{25'd667924}}, '{'{25'd0}}, '{'{25'd190836}}, '{'{25'd1288140}}, '{'{-25'd1526684}}},
    '{'{'{-25'd1560016}}, '{'{-25'd288892}}, '{'{-25'd1675573}}, '{'{25'd1733351}}, '{'{25'd1271124}}, '{'{-25'd288892}}, '{'{25'd7337854}}, '{'{-25'd635562}}, '{'{25'd346670}}, '{'{25'd3640038}}, '{'{-25'd1502238}}, '{'{25'd1848908}}, '{'{25'd1502238}}, '{'{-25'd1906687}}, '{'{-25'd1097789}}, '{'{25'd693341}}, '{'{-25'd2080022}}, '{'{-25'd866676}}, '{'{25'd231114}}, '{'{-25'd3120033}}, '{'{25'd4275600}}, '{'{-25'd982232}}, '{'{25'd1848908}}, '{'{-25'd1097789}}, '{'{-25'd1040011}}, '{'{-25'd1097789}}, '{'{-25'd924454}}, '{'{25'd577784}}, '{'{25'd1328903}}, '{'{25'd2888919}}, '{'{-25'd577784}}, '{'{25'd2137800}}, '{'{-25'd751119}}, '{'{-25'd1560016}}, '{'{25'd1791130}}, '{'{-25'd808897}}, '{'{-25'd2080022}}, '{'{-25'd924454}}, '{'{25'd1906687}}, '{'{25'd1271124}}, '{'{-25'd3235589}}, '{'{25'd346670}}, '{'{-25'd1617795}}, '{'{-25'd1444460}}, '{'{-25'd751119}}, '{'{-25'd808897}}, '{'{25'd1097789}}, '{'{-25'd1560016}}, '{'{25'd1848908}}, '{'{25'd1675573}}, '{'{25'd2484470}}, '{'{-25'd1213346}}, '{'{25'd751119}}, '{'{-25'd288892}}, '{'{25'd2773362}}, '{'{-25'd462227}}, '{'{-25'd1560016}}, '{'{-25'd462227}}, '{'{-25'd1617795}}, '{'{-25'd231114}}, '{'{25'd924454}}, '{'{25'd5026719}}, '{'{-25'd1097789}}, '{'{-25'd635562}}},
    '{'{'{25'd469723}}, '{'{-25'd858921}}, '{'{25'd993128}}, '{'{-25'd778398}}, '{'{25'd805239}}, '{'{25'd228151}}, '{'{25'd1409168}}, '{'{25'd496564}}, '{'{-25'd885763}}, '{'{25'd147627}}, '{'{-25'd228151}}, '{'{-25'd1704422}}, '{'{25'd590508}}, '{'{-25'd1637319}}, '{'{-25'd1382327}}, '{'{-25'd335516}}, '{'{-25'd1140755}}, '{'{25'd214730}}, '{'{25'd1248120}}, '{'{25'd1248120}}, '{'{-25'd1382327}}, '{'{25'd13421}}, '{'{-25'd912604}}, '{'{25'd1342065}}, '{'{-25'd1288382}}, '{'{-25'd872342}}, '{'{-25'd1248120}}, '{'{-25'd1181017}}, '{'{25'd1087072}}, '{'{25'd1181017}}, '{'{-25'd845501}}, '{'{-25'd174468}}, '{'{25'd120786}}, '{'{25'd483143}}, '{'{-25'd617350}}, '{'{-25'd603929}}, '{'{25'd1127334}}, '{'{25'd134206}}, '{'{25'd93945}}, '{'{-25'd1691002}}, '{'{-25'd536826}}, '{'{25'd751556}}, '{'{25'd845501}}, '{'{-25'd1409168}}, '{'{-25'd1033390}}, '{'{-25'd1060231}}, '{'{25'd1234700}}, '{'{-25'd1087072}}, '{'{-25'd93945}}, '{'{25'd469723}}, '{'{25'd1462851}}, '{'{-25'd362357}}, '{'{-25'd939445}}, '{'{-25'd107365}}, '{'{25'd1046811}}, '{'{25'd1113914}}, '{'{-25'd214730}}, '{'{-25'd1181017}}, '{'{-25'd1006549}}, '{'{-25'd751556}}, '{'{-25'd657612}}, '{'{-25'd603929}}, '{'{25'd1476271}}, '{'{-25'd469723}}},
    '{'{'{-25'd837381}}, '{'{25'd942054}}, '{'{-25'd1116508}}, '{'{25'd488472}}, '{'{25'd1151399}}, '{'{-25'd523363}}, '{'{-25'd17445}}, '{'{25'd0}}, '{'{25'd1221181}}, '{'{-25'd662927}}, '{'{25'd1727099}}, '{'{25'd1639871}}, '{'{25'd645481}}, '{'{25'd1744544}}, '{'{25'd523363}}, '{'{25'd348909}}, '{'{-25'd819936}}, '{'{25'd1081617}}, '{'{-25'd1064172}}, '{'{-25'd1343299}}, '{'{-25'd2128344}}, '{'{25'd1116508}}, '{'{25'd1186290}}, '{'{25'd732709}}, '{'{-25'd1011836}}, '{'{-25'd662927}}, '{'{25'd750154}}, '{'{-25'd1552644}}, '{'{25'd540809}}, '{'{-25'd976945}}, '{'{25'd261682}}, '{'{-25'd1360744}}, '{'{25'd1692208}}, '{'{-25'd1029281}}, '{'{25'd1570090}}, '{'{25'd942054}}, '{'{-25'd540809}}, '{'{-25'd17445}}, '{'{-25'd1482862}}, '{'{-25'd959499}}, '{'{-25'd1849217}}, '{'{25'd1465417}}, '{'{-25'd1517753}}, '{'{25'd907163}}, '{'{25'd837381}}, '{'{25'd1779435}}, '{'{25'd1587535}}, '{'{25'd1744544}}, '{'{25'd139564}}, '{'{-25'd1011836}}, '{'{25'd1186290}}, '{'{-25'd662927}}, '{'{-25'd1500308}}, '{'{-25'd436136}}, '{'{25'd69782}}, '{'{25'd662927}}, '{'{25'd1203735}}, '{'{25'd715263}}, '{'{-25'd2215571}}, '{'{25'd1064172}}, '{'{-25'd610590}}, '{'{-25'd1692208}}, '{'{-25'd1413081}}, '{'{-25'd785045}}},
    '{'{'{-25'd1070021}}, '{'{25'd189842}}, '{'{25'd1674066}}, '{'{25'd396943}}, '{'{-25'd1190830}}, '{'{25'd1018246}}, '{'{25'd224359}}, '{'{-25'd396943}}, '{'{-25'd327910}}, '{'{-25'd310651}}, '{'{25'd1656807}}, '{'{25'd1208089}}, '{'{25'd1380673}}, '{'{25'd17258}}, '{'{-25'd17258}}, '{'{25'd362427}}, '{'{-25'd1639549}}, '{'{-25'd1156313}}, '{'{-25'd1225347}}, '{'{-25'd983729}}, '{'{25'd1984717}}, '{'{-25'd897437}}, '{'{25'd862920}}, '{'{-25'd1242605}}, '{'{-25'd327910}}, '{'{-25'd1070021}}, '{'{-25'd414202}}, '{'{25'd1000988}}, '{'{25'd742112}}, '{'{25'd655819}}, '{'{25'd1070021}}, '{'{25'd1898425}}, '{'{25'd1518740}}, '{'{25'd1070021}}, '{'{25'd845662}}, '{'{25'd1277122}}, '{'{-25'd1466965}}, '{'{25'd448719}}, '{'{25'd2191818}}, '{'{25'd86292}}, '{'{25'd241618}}, '{'{25'd1622290}}, '{'{25'd500494}}, '{'{25'd1725841}}, '{'{-25'd310651}}, '{'{-25'd1208089}}, '{'{25'd1553257}}, '{'{-25'd1277122}}, '{'{25'd155326}}, '{'{-25'd17258}}, '{'{-25'd1432448}}, '{'{25'd983729}}, '{'{25'd1225347}}, '{'{-25'd793887}}, '{'{25'd1104538}}, '{'{25'd258876}}, '{'{-25'd1656807}}, '{'{25'd345168}}, '{'{25'd845662}}, '{'{-25'd362427}}, '{'{-25'd431460}}, '{'{-25'd1156313}}, '{'{25'd811145}}, '{'{-25'd138067}}},
    '{'{'{-25'd1656603}}, '{'{-25'd1411714}}, '{'{-25'd14405}}, '{'{25'd1094798}}, '{'{25'd864314}}, '{'{-25'd1094798}}, '{'{25'd950746}}, '{'{-25'd878720}}, '{'{25'd677046}}, '{'{25'd1195635}}, '{'{25'd460968}}, '{'{25'd1498145}}, '{'{-25'd1080393}}, '{'{-25'd1843871}}, '{'{-25'd648236}}, '{'{25'd1397308}}, '{'{25'd1282066}}, '{'{-25'd1152419}}, '{'{-25'd374536}}, '{'{-25'd532994}}, '{'{25'd835504}}, '{'{25'd777883}}, '{'{-25'd1843871}}, '{'{-25'd86431}}, '{'{-25'd475373}}, '{'{25'd864314}}, '{'{-25'd302510}}, '{'{-25'd388941}}, '{'{25'd187268}}, '{'{-25'd244889}}, '{'{-25'd1080393}}, '{'{25'd1123609}}, '{'{25'd504183}}, '{'{25'd14405}}, '{'{-25'd1065988}}, '{'{-25'd1282066}}, '{'{25'd0}}, '{'{-25'd1642197}}, '{'{-25'd72026}}, '{'{-25'd936341}}, '{'{25'd1829465}}, '{'{-25'd1440524}}, '{'{25'd1714224}}, '{'{-25'd1310877}}, '{'{-25'd1238851}}, '{'{25'd561804}}, '{'{25'd446562}}, '{'{25'd1699818}}, '{'{25'd936341}}, '{'{-25'd1296472}}, '{'{-25'd57621}}, '{'{25'd1829465}}, '{'{25'd1037177}}, '{'{25'd288105}}, '{'{25'd331321}}, '{'{-25'd576210}}, '{'{25'd1181230}}, '{'{25'd1671008}}, '{'{-25'd1685413}}, '{'{25'd259294}}, '{'{25'd1368498}}, '{'{25'd1786250}}, '{'{25'd1526955}}, '{'{25'd1210040}}},
    '{'{'{25'd1259106}}, '{'{25'd2064933}}, '{'{-25'd1007284}}, '{'{-25'd302185}}, '{'{25'd654735}}, '{'{25'd50364}}, '{'{25'd5892614}}, '{'{-25'd1561291}}, '{'{25'd705099}}, '{'{-25'd6446621}}, '{'{25'd1712384}}, '{'{25'd705099}}, '{'{-25'd1259106}}, '{'{-25'd3525496}}, '{'{-25'd805828}}, '{'{25'd856192}}, '{'{25'd1057649}}, '{'{-25'd906556}}, '{'{-25'd2367118}}, '{'{25'd755463}}, '{'{25'd0}}, '{'{-25'd604371}}, '{'{-25'd201457}}, '{'{-25'd1662019}}, '{'{-25'd755463}}, '{'{25'd1108013}}, '{'{25'd100728}}, '{'{-25'd1007284}}, '{'{25'd151093}}, '{'{25'd1964205}}, '{'{25'd2921125}}, '{'{25'd1913840}}, '{'{-25'd1662019}}, '{'{25'd352550}}, '{'{-25'd302185}}, '{'{-25'd1108013}}, '{'{-25'd1108013}}, '{'{25'd604371}}, '{'{25'd2820397}}, '{'{-25'd1561291}}, '{'{-25'd3273675}}, '{'{25'd705099}}, '{'{-25'd2216026}}, '{'{25'd1158377}}, '{'{-25'd1611655}}, '{'{25'd1158377}}, '{'{-25'd1108013}}, '{'{-25'd956920}}, '{'{-25'd956920}}, '{'{25'd1208741}}, '{'{25'd2568575}}, '{'{-25'd1309470}}, '{'{-25'd352550}}, '{'{25'd1359834}}, '{'{25'd2115297}}, '{'{25'd453278}}, '{'{-25'd1561291}}, '{'{-25'd251821}}, '{'{25'd201457}}, '{'{25'd201457}}, '{'{-25'd1510927}}, '{'{25'd4583144}}, '{'{-25'd1359834}}, '{'{25'd1158377}}},
    '{'{'{-25'd764752}}, '{'{25'd224927}}, '{'{-25'd794742}}, '{'{25'd1574489}}, '{'{-25'd1229601}}, '{'{-25'd644791}}, '{'{25'd1724440}}, '{'{-25'd74976}}, '{'{-25'd1664460}}, '{'{-25'd1094645}}, '{'{25'd1544499}}, '{'{-25'd884713}}, '{'{-25'd344888}}, '{'{25'd479844}}, '{'{25'd494839}}, '{'{25'd614800}}, '{'{25'd509834}}, '{'{-25'd764752}}, '{'{25'd674781}}, '{'{25'd1409542}}, '{'{25'd239922}}, '{'{25'd1064654}}, '{'{-25'd674781}}, '{'{25'd764752}}, '{'{25'd509834}}, '{'{25'd164946}}, '{'{25'd1364557}}, '{'{25'd1784421}}, '{'{-25'd599805}}, '{'{-25'd1799416}}, '{'{25'd749757}}, '{'{25'd1034664}}, '{'{25'd1514508}}, '{'{25'd629796}}, '{'{25'd119961}}, '{'{-25'd494839}}, '{'{25'd1034664}}, '{'{-25'd1124635}}, '{'{25'd1079649}}, '{'{-25'd1904382}}, '{'{25'd1709445}}, '{'{25'd194937}}, '{'{-25'd1589484}}, '{'{25'd389873}}, '{'{25'd1229601}}, '{'{25'd1184615}}, '{'{25'd1379552}}, '{'{-25'd104966}}, '{'{25'd1499513}}, '{'{25'd614800}}, '{'{25'd1514508}}, '{'{25'd1694450}}, '{'{25'd209932}}, '{'{-25'd1274586}}, '{'{25'd74976}}, '{'{-25'd794742}}, '{'{-25'd194937}}, '{'{-25'd239922}}, '{'{25'd284908}}, '{'{-25'd704771}}, '{'{25'd1424538}}, '{'{25'd1334567}}, '{'{25'd1244596}}, '{'{25'd329893}}},
    '{'{'{25'd1319226}}, '{'{25'd253185}}, '{'{25'd1319226}}, '{'{-25'd519695}}, '{'{25'd413091}}, '{'{25'd652950}}, '{'{25'd26651}}, '{'{-25'd1465807}}, '{'{25'd133255}}, '{'{25'd1106018}}, '{'{-25'd932786}}, '{'{-25'd159906}}, '{'{25'd133255}}, '{'{25'd666276}}, '{'{25'd1212622}}, '{'{-25'd812857}}, '{'{-25'd319812}}, '{'{-25'd1492458}}, '{'{-25'd1066041}}, '{'{25'd1599062}}, '{'{25'd1199297}}, '{'{25'd1225948}}, '{'{-25'd1705666}}, '{'{25'd1399179}}, '{'{25'd1412505}}, '{'{-25'd599648}}, '{'{25'd1585737}}, '{'{-25'd159906}}, '{'{25'd479719}}, '{'{25'd1145994}}, '{'{-25'd572997}}, '{'{25'd479719}}, '{'{-25'd359789}}, '{'{-25'd119930}}, '{'{-25'd1012739}}, '{'{-25'd1039390}}, '{'{25'd1372528}}, '{'{-25'd13326}}, '{'{-25'd1505783}}, '{'{-25'd999414}}, '{'{25'd759554}}, '{'{-25'd1012739}}, '{'{25'd133255}}, '{'{-25'd1599062}}, '{'{-25'd79953}}, '{'{-25'd1145994}}, '{'{-25'd133255}}, '{'{-25'd919461}}, '{'{-25'd1625713}}, '{'{-25'd972763}}, '{'{-25'd533021}}, '{'{25'd1519109}}, '{'{-25'd786206}}, '{'{-25'd1052716}}, '{'{-25'd253185}}, '{'{-25'd1399179}}, '{'{25'd39977}}, '{'{25'd26651}}, '{'{-25'd1185971}}, '{'{25'd932786}}, '{'{25'd692927}}, '{'{-25'd293161}}, '{'{25'd1532434}}, '{'{25'd1145994}}},
    '{'{'{-25'd1315404}}, '{'{-25'd575489}}, '{'{25'd295966}}, '{'{-25'd1068766}}, '{'{-25'd1644255}}, '{'{-25'd197311}}, '{'{25'd1594927}}, '{'{25'd1216749}}, '{'{25'd756357}}, '{'{25'd1710025}}, '{'{25'd1019438}}, '{'{-25'd1150979}}, '{'{25'd1150979}}, '{'{-25'd1858008}}, '{'{25'd1183864}}, '{'{-25'd295966}}, '{'{25'd411064}}, '{'{25'd739915}}, '{'{25'd312408}}, '{'{25'd509719}}, '{'{25'd476834}}, '{'{25'd230196}}, '{'{25'd1019438}}, '{'{25'd1545600}}, '{'{25'd427506}}, '{'{25'd230196}}, '{'{-25'd789242}}, '{'{25'd707030}}, '{'{25'd147983}}, '{'{25'd394621}}, '{'{-25'd1052323}}, '{'{-25'd312408}}, '{'{25'd542604}}, '{'{25'd180868}}, '{'{25'd1052323}}, '{'{-25'd1512715}}, '{'{-25'd937225}}, '{'{-25'd98655}}, '{'{-25'd1068766}}, '{'{25'd16443}}, '{'{25'd1496272}}, '{'{-25'd559047}}, '{'{25'd460391}}, '{'{25'd1463387}}, '{'{-25'd953668}}, '{'{-25'd82213}}, '{'{25'd82213}}, '{'{25'd1381174}}, '{'{-25'd197311}}, '{'{-25'd855013}}, '{'{-25'd937225}}, '{'{-25'd2104647}}, '{'{25'd49328}}, '{'{-25'd1381174}}, '{'{-25'd2088204}}, '{'{25'd1019438}}, '{'{-25'd542604}}, '{'{25'd1611370}}, '{'{-25'd164426}}, '{'{-25'd1315404}}, '{'{-25'd1529157}}, '{'{-25'd1019438}}, '{'{-25'd1085208}}, '{'{25'd575489}}},
    '{'{'{-25'd274328}}, '{'{25'd2011737}}, '{'{25'd274328}}, '{'{-25'd1554524}}, '{'{-25'd1645966}}, '{'{25'd1097311}}, '{'{25'd1005868}}, '{'{25'd640098}}, '{'{25'd457213}}, '{'{25'd7223963}}, '{'{-25'd365770}}, '{'{-25'd731541}}, '{'{25'd1280196}}, '{'{25'd1371639}}, '{'{25'd731541}}, '{'{-25'd1188753}}, '{'{25'd0}}, '{'{-25'd548655}}, '{'{25'd1828851}}, '{'{-25'd4206358}}, '{'{25'd1005868}}, '{'{25'd1737409}}, '{'{25'd457213}}, '{'{-25'd1463081}}, '{'{-25'd640098}}, '{'{-25'd457213}}, '{'{-25'd1828851}}, '{'{25'd1097311}}, '{'{-25'd365770}}, '{'{25'd2011737}}, '{'{25'd2834720}}, '{'{25'd1188753}}, '{'{25'd3840588}}, '{'{-25'd1737409}}, '{'{-25'd1280196}}, '{'{25'd2011737}}, '{'{25'd1645966}}, '{'{25'd548655}}, '{'{-25'd3291933}}, '{'{25'd3200490}}, '{'{-25'd1920294}}, '{'{25'd1645966}}, '{'{-25'd1737409}}, '{'{25'd1280196}}, '{'{25'd1280196}}, '{'{-25'd274328}}, '{'{-25'd1280196}}, '{'{25'd91443}}, '{'{25'd457213}}, '{'{25'd548655}}, '{'{-25'd6675308}}, '{'{25'd274328}}, '{'{-25'd822983}}, '{'{-25'd822983}}, '{'{25'd1280196}}, '{'{-25'd1463081}}, '{'{-25'd274328}}, '{'{-25'd1371639}}, '{'{-25'd1645966}}, '{'{25'd274328}}, '{'{25'd731541}}, '{'{25'd11613206}}, '{'{-25'd1005868}}, '{'{25'd182885}}},
    '{'{'{25'd245997}}, '{'{25'd1632528}}, '{'{25'd290724}}, '{'{25'd335451}}, '{'{25'd849809}}, '{'{25'd1364167}}, '{'{25'd201271}}, '{'{-25'd760355}}, '{'{-25'd1073443}}, '{'{25'd805082}}, '{'{-25'd156544}}, '{'{25'd447268}}, '{'{-25'd1319440}}, '{'{-25'd156544}}, '{'{-25'd939263}}, '{'{25'd760355}}, '{'{-25'd313088}}, '{'{25'd514358}}, '{'{25'd1453621}}, '{'{25'd1364167}}, '{'{25'd2840151}}, '{'{-25'd380178}}, '{'{-25'd201271}}, '{'{25'd894536}}, '{'{-25'd1252350}}, '{'{25'd424905}}, '{'{25'd827446}}, '{'{-25'd1386531}}, '{'{25'd1677255}}, '{'{25'd782719}}, '{'{25'd22363}}, '{'{25'd715629}}, '{'{25'd1453621}}, '{'{25'd1475984}}, '{'{-25'd1118170}}, '{'{25'd0}}, '{'{-25'd827446}}, '{'{-25'd89454}}, '{'{25'd268361}}, '{'{-25'd715629}}, '{'{25'd424905}}, '{'{-25'd1207623}}, '{'{25'd1408894}}, '{'{25'd1051080}}, '{'{-25'd693265}}, '{'{-25'd491995}}, '{'{25'd1207623}}, '{'{25'd1118170}}, '{'{25'd357814}}, '{'{25'd1028716}}, '{'{25'd983989}}, '{'{-25'd1386531}}, '{'{-25'd1341804}}, '{'{-25'd1520711}}, '{'{25'd1520711}}, '{'{-25'd983989}}, '{'{25'd760355}}, '{'{-25'd1632528}}, '{'{25'd111817}}, '{'{-25'd827446}}, '{'{25'd178907}}, '{'{25'd939263}}, '{'{25'd827446}}, '{'{25'd268361}}},
    '{'{'{25'd532182}}, '{'{-25'd177394}}, '{'{25'd1655677}}, '{'{-25'd1064364}}, '{'{25'd1360020}}, '{'{-25'd236525}}, '{'{-25'd295657}}, '{'{-25'd1123495}}, '{'{25'd1478283}}, '{'{-25'd1005232}}, '{'{-25'd1182626}}, '{'{25'd1123495}}, '{'{-25'd177394}}, '{'{25'd532182}}, '{'{-25'd650444}}, '{'{25'd118263}}, '{'{25'd1773939}}, '{'{25'd1360020}}, '{'{-25'd118263}}, '{'{25'd1005232}}, '{'{25'd3725273}}, '{'{25'd1064364}}, '{'{-25'd236525}}, '{'{-25'd1005232}}, '{'{25'd1596545}}, '{'{-25'd1182626}}, '{'{-25'd1478283}}, '{'{-25'd1478283}}, '{'{-25'd1360020}}, '{'{25'd2838303}}, '{'{25'd1714808}}, '{'{-25'd177394}}, '{'{25'd2601778}}, '{'{-25'd177394}}, '{'{-25'd827838}}, '{'{25'd886970}}, '{'{-25'd946101}}, '{'{-25'd1300889}}, '{'{-25'd1182626}}, '{'{25'd236525}}, '{'{25'd7509676}}, '{'{25'd1005232}}, '{'{-25'd177394}}, '{'{-25'd532182}}, '{'{25'd295657}}, '{'{25'd59131}}, '{'{-25'd59131}}, '{'{25'd1064364}}, '{'{-25'd1123495}}, '{'{25'd236525}}, '{'{-25'd2424384}}, '{'{25'd295657}}, '{'{-25'd118263}}, '{'{-25'd1596545}}, '{'{-25'd768707}}, '{'{-25'd768707}}, '{'{25'd768707}}, '{'{-25'd236525}}, '{'{25'd1478283}}, '{'{25'd1419151}}, '{'{25'd946101}}, '{'{25'd473050}}, '{'{25'd886970}}, '{'{-25'd946101}}},
    '{'{'{25'd1372862}}, '{'{25'd964714}}, '{'{25'd1632593}}, '{'{-25'd1113131}}, '{'{25'd1298653}}, '{'{-25'd779192}}, '{'{25'd1001818}}, '{'{25'd445253}}, '{'{25'd1261549}}, '{'{25'd259731}}, '{'{-25'd704983}}, '{'{-25'd1558384}}, '{'{-25'd519461}}, '{'{-25'd742088}}, '{'{25'd556566}}, '{'{-25'd111313}}, '{'{25'd816296}}, '{'{-25'd1632593}}, '{'{25'd1781010}}, '{'{-25'd1929428}}, '{'{25'd4712256}}, '{'{25'd927609}}, '{'{25'd779192}}, '{'{25'd1076027}}, '{'{-25'd1224444}}, '{'{25'd259731}}, '{'{25'd1335758}}, '{'{-25'd74209}}, '{'{25'd704983}}, '{'{-25'd185522}}, '{'{-25'd37104}}, '{'{-25'd482357}}, '{'{25'd964714}}, '{'{-25'd222626}}, '{'{-25'd259731}}, '{'{25'd111313}}, '{'{25'd222626}}, '{'{-25'd1113131}}, '{'{25'd593670}}, '{'{-25'd1298653}}, '{'{-25'd1781010}}, '{'{-25'd1113131}}, '{'{25'd1113131}}, '{'{25'd1632593}}, '{'{25'd185522}}, '{'{25'd853401}}, '{'{-25'd1076027}}, '{'{25'd1706801}}, '{'{25'd519461}}, '{'{25'd964714}}, '{'{-25'd779192}}, '{'{25'd704983}}, '{'{-25'd1261549}}, '{'{25'd1595488}}, '{'{-25'd1335758}}, '{'{-25'd779192}}, '{'{25'd1447071}}, '{'{25'd1372862}}, '{'{-25'd593670}}, '{'{25'd1150236}}, '{'{-25'd1521279}}, '{'{-25'd2263367}}, '{'{-25'd1038923}}, '{'{-25'd630774}}},
    '{'{'{25'd1328685}}, '{'{-25'd47453}}, '{'{25'd31635}}, '{'{25'd2008845}}, '{'{-25'd142359}}, '{'{25'd1597585}}, '{'{-25'd695978}}, '{'{25'd363806}}, '{'{-25'd173994}}, '{'{25'd996513}}, '{'{-25'd253083}}, '{'{25'd1328685}}, '{'{-25'd1407773}}, '{'{-25'd806701}}, '{'{-25'd506166}}, '{'{25'd1407773}}, '{'{-25'd1771579}}, '{'{25'd1328685}}, '{'{-25'd743431}}, '{'{25'd458713}}, '{'{25'd458713}}, '{'{25'd1439408}}, '{'{-25'd711795}}, '{'{-25'd221447}}, '{'{25'd1629220}}, '{'{-25'd158177}}, '{'{25'd1154690}}, '{'{25'd79088}}, '{'{25'd1502679}}, '{'{-25'd759248}}, '{'{-25'd664342}}, '{'{-25'd980696}}, '{'{-25'd173994}}, '{'{25'd1281232}}, '{'{25'd47453}}, '{'{25'd1217961}}, '{'{-25'd284718}}, '{'{25'd1518497}}, '{'{25'd1882303}}, '{'{25'd933243}}, '{'{-25'd616889}}, '{'{25'd743431}}, '{'{-25'd980696}}, '{'{-25'd711795}}, '{'{-25'd1012331}}, '{'{25'd1059784}}, '{'{-25'd411260}}, '{'{25'd1502679}}, '{'{25'd1581767}}, '{'{25'd1107237}}, '{'{25'd1423591}}, '{'{25'd442895}}, '{'{25'd1645038}}, '{'{-25'd1186326}}, '{'{25'd1597585}}, '{'{-25'd15818}}, '{'{25'd1407773}}, '{'{25'd379624}}, '{'{-25'd63271}}, '{'{-25'd1281232}}, '{'{-25'd680160}}, '{'{25'd47453}}, '{'{25'd996513}}, '{'{25'd1423591}}},
    '{'{'{25'd18671}}, '{'{-25'd784166}}, '{'{25'd1605674}}, '{'{-25'd1474980}}, '{'{-25'd1026885}}, '{'{25'd112024}}, '{'{-25'd1400297}}, '{'{25'd989543}}, '{'{-25'd149365}}, '{'{25'd2016428}}, '{'{25'd429424}}, '{'{-25'd634801}}, '{'{25'd709484}}, '{'{25'd2371170}}, '{'{25'd1624345}}, '{'{25'd1643015}}, '{'{25'd1250932}}, '{'{-25'd1306944}}, '{'{-25'd802837}}, '{'{-25'd373413}}, '{'{25'd2371170}}, '{'{25'd653472}}, '{'{-25'd298730}}, '{'{-25'd933531}}, '{'{-25'd1418968}}, '{'{-25'd765496}}, '{'{25'd1418968}}, '{'{-25'd877520}}, '{'{25'd634801}}, '{'{25'd1288273}}, '{'{-25'd373413}}, '{'{25'd354742}}, '{'{-25'd448095}}, '{'{25'd1026885}}, '{'{25'd392083}}, '{'{-25'd1680357}}, '{'{-25'd1587003}}, '{'{25'd1250932}}, '{'{25'd2240475}}, '{'{-25'd672143}}, '{'{-25'd541448}}, '{'{-25'd1568333}}, '{'{-25'd821508}}, '{'{-25'd728154}}, '{'{25'd373413}}, '{'{25'd1512321}}, '{'{-25'd858849}}, '{'{25'd728154}}, '{'{-25'd840178}}, '{'{-25'd522778}}, '{'{25'd466766}}, '{'{-25'd840178}}, '{'{25'd1194920}}, '{'{25'd672143}}, '{'{25'd1568333}}, '{'{-25'd802837}}, '{'{25'd1344285}}, '{'{-25'd952202}}, '{'{25'd466766}}, '{'{25'd1530991}}, '{'{-25'd728154}}, '{'{-25'd1269603}}, '{'{25'd578789}}, '{'{25'd186706}}},
    '{'{'{-25'd1552781}}, '{'{25'd221826}}, '{'{-25'd369710}}, '{'{25'd739420}}, '{'{-25'd1404897}}, '{'{25'd1552781}}, '{'{25'd9390630}}, '{'{25'd591536}}, '{'{25'd665478}}, '{'{25'd5619590}}, '{'{-25'd591536}}, '{'{-25'd1626723}}, '{'{25'd1478839}}, '{'{25'd2735853}}, '{'{25'd887304}}, '{'{25'd961246}}, '{'{-25'd1035188}}, '{'{-25'd295768}}, '{'{25'd0}}, '{'{25'd665478}}, '{'{25'd4214692}}, '{'{-25'd665478}}, '{'{25'd3031621}}, '{'{-25'd1626723}}, '{'{25'd295768}}, '{'{-25'd961246}}, '{'{25'd887304}}, '{'{25'd2587969}}, '{'{25'd1257013}}, '{'{25'd739420}}, '{'{-25'd591536}}, '{'{25'd1700665}}, '{'{25'd73942}}, '{'{-25'd517594}}, '{'{25'd1478839}}, '{'{25'd221826}}, '{'{-25'd1035188}}, '{'{-25'd517594}}, '{'{-25'd517594}}, '{'{25'd1109130}}, '{'{-25'd6950545}}, '{'{-25'd1404897}}, '{'{-25'd2218259}}, '{'{25'd369710}}, '{'{25'd961246}}, '{'{-25'd443652}}, '{'{25'd1478839}}, '{'{25'd1552781}}, '{'{25'd369710}}, '{'{-25'd1404897}}, '{'{-25'd2218259}}, '{'{-25'd3844982}}, '{'{-25'd2144317}}, '{'{-25'd2144317}}, '{'{25'd1848549}}, '{'{25'd1700665}}, '{'{25'd813362}}, '{'{-25'd887304}}, '{'{25'd1404897}}, '{'{25'd1552781}}, '{'{-25'd1552781}}, '{'{-25'd591536}}, '{'{25'd1774607}}, '{'{-25'd443652}}},
    '{'{'{25'd504503}}, '{'{25'd917277}}, '{'{25'd458639}}, '{'{25'd2981152}}, '{'{25'd91728}}, '{'{25'd1559372}}, '{'{-25'd5870575}}, '{'{25'd963141}}, '{'{25'd366911}}, '{'{-25'd2247330}}, '{'{-25'd504503}}, '{'{25'd504503}}, '{'{25'd137592}}, '{'{-25'd2476649}}, '{'{-25'd825550}}, '{'{25'd1742827}}, '{'{25'd458639}}, '{'{-25'd458639}}, '{'{-25'd321047}}, '{'{-25'd1880419}}, '{'{-25'd5090890}}, '{'{-25'd504503}}, '{'{25'd366911}}, '{'{25'd137592}}, '{'{25'd1100733}}, '{'{-25'd687958}}, '{'{25'd779686}}, '{'{25'd366911}}, '{'{25'd550366}}, '{'{25'd4861570}}, '{'{-25'd1559372}}, '{'{25'd642094}}, '{'{25'd1009005}}, '{'{-25'd1605235}}, '{'{-25'd1421780}}, '{'{-25'd412775}}, '{'{25'd1467644}}, '{'{-25'd871414}}, '{'{25'd1100733}}, '{'{-25'd733822}}, '{'{-25'd1330052}}, '{'{25'd1192461}}, '{'{-25'd1742827}}, '{'{-25'd458639}}, '{'{25'd1605235}}, '{'{-25'd45864}}, '{'{25'd504503}}, '{'{-25'd275183}}, '{'{-25'd825550}}, '{'{25'd229319}}, '{'{25'd321047}}, '{'{25'd1696963}}, '{'{-25'd45864}}, '{'{-25'd687958}}, '{'{25'd1880419}}, '{'{25'd1330052}}, '{'{25'd550366}}, '{'{-25'd1421780}}, '{'{-25'd1238324}}, '{'{25'd687958}}, '{'{25'd458639}}, '{'{25'd4402932}}, '{'{-25'd917277}}, '{'{-25'd183455}}},
    '{'{'{25'd1582835}}, '{'{25'd1074585}}, '{'{-25'd726071}}, '{'{25'd1452142}}, '{'{25'd871285}}, '{'{25'd1306928}}, '{'{25'd842243}}, '{'{25'd1481185}}, '{'{25'd377557}}, '{'{25'd726071}}, '{'{-25'd1553792}}, '{'{-25'd1684485}}, '{'{-25'd697028}}, '{'{-25'd537293}}, '{'{-25'd1335971}}, '{'{-25'd842243}}, '{'{25'd1466664}}, '{'{-25'd261386}}, '{'{25'd493728}}, '{'{25'd392078}}, '{'{25'd769636}}, '{'{25'd1423100}}, '{'{-25'd377557}}, '{'{-25'd290428}}, '{'{25'd58086}}, '{'{25'd943893}}, '{'{25'd464686}}, '{'{-25'd740593}}, '{'{25'd319471}}, '{'{-25'd522771}}, '{'{-25'd1553792}}, '{'{-25'd508250}}, '{'{25'd1786135}}, '{'{25'd711550}}, '{'{25'd1031021}}, '{'{-25'd1423100}}, '{'{-25'd1452142}}, '{'{25'd101650}}, '{'{-25'd697028}}, '{'{25'd1844221}}, '{'{25'd827721}}, '{'{25'd1219800}}, '{'{25'd595378}}, '{'{-25'd1335971}}, '{'{25'd1001978}}, '{'{25'd871285}}, '{'{-25'd972935}}, '{'{25'd1699007}}, '{'{25'd1031021}}, '{'{25'd1394057}}, '{'{25'd14521}}, '{'{-25'd1103628}}, '{'{25'd159736}}, '{'{25'd464686}}, '{'{25'd1292407}}, '{'{25'd624421}}, '{'{-25'd464686}}, '{'{-25'd798678}}, '{'{-25'd900328}}, '{'{25'd217821}}, '{'{25'd711550}}, '{'{-25'd1016500}}, '{'{25'd1452142}}, '{'{-25'd464686}}},
    '{'{'{25'd649674}}, '{'{-25'd949524}}, '{'{-25'd649674}}, '{'{25'd249875}}, '{'{-25'd1449273}}, '{'{25'd699649}}, '{'{25'd2248873}}, '{'{25'd1699148}}, '{'{-25'd999499}}, '{'{-25'd3348321}}, '{'{25'd699649}}, '{'{25'd599699}}, '{'{-25'd1549223}}, '{'{-25'd649674}}, '{'{25'd199900}}, '{'{25'd1599198}}, '{'{-25'd899549}}, '{'{25'd1699148}}, '{'{-25'd1249374}}, '{'{25'd2298848}}, '{'{-25'd6346818}}, '{'{-25'd1649173}}, '{'{25'd999499}}, '{'{-25'd1099449}}, '{'{-25'd1299349}}, '{'{25'd999499}}, '{'{-25'd1049474}}, '{'{25'd1099449}}, '{'{-25'd749624}}, '{'{25'd1849073}}, '{'{-25'd449775}}, '{'{25'd1099449}}, '{'{-25'd199900}}, '{'{25'd599699}}, '{'{25'd299850}}, '{'{-25'd1549223}}, '{'{25'd299850}}, '{'{-25'd749624}}, '{'{25'd499749}}, '{'{-25'd249875}}, '{'{-25'd3098447}}, '{'{25'd2148923}}, '{'{-25'd449775}}, '{'{-25'd499749}}, '{'{25'd349825}}, '{'{-25'd449775}}, '{'{-25'd1699148}}, '{'{-25'd1199399}}, '{'{-25'd1149424}}, '{'{-25'd49975}}, '{'{25'd449775}}, '{'{-25'd849574}}, '{'{25'd399800}}, '{'{25'd1099449}}, '{'{25'd1149424}}, '{'{25'd1599198}}, '{'{-25'd1649173}}, '{'{25'd1049474}}, '{'{25'd1249374}}, '{'{25'd699649}}, '{'{25'd1449273}}, '{'{25'd2498747}}, '{'{-25'd399800}}, '{'{-25'd1299349}}},
    '{'{'{25'd491894}}, '{'{-25'd532885}}, '{'{25'd1339045}}, '{'{-25'd286938}}, '{'{-25'd54655}}, '{'{25'd970124}}, '{'{-25'd1120425}}, '{'{-25'd1175080}}, '{'{25'd942797}}, '{'{-25'd27327}}, '{'{-25'd95646}}, '{'{-25'd1243399}}, '{'{25'd1175080}}, '{'{-25'd1311717}}, '{'{-25'd573876}}, '{'{-25'd1038443}}, '{'{-25'd382584}}, '{'{-25'd765168}}, '{'{25'd888142}}, '{'{25'd273274}}, '{'{25'd956461}}, '{'{25'd1216071}}, '{'{25'd1161416}}, '{'{-25'd245947}}, '{'{25'd1011115}}, '{'{25'd724177}}, '{'{-25'd478230}}, '{'{25'd13664}}, '{'{-25'd1434691}}, '{'{-25'd765168}}, '{'{25'd204956}}, '{'{25'd1571328}}, '{'{-25'd491894}}, '{'{-25'd95646}}, '{'{-25'd860815}}, '{'{25'd505558}}, '{'{-25'd1735293}}, '{'{25'd519221}}, '{'{-25'd1270726}}, '{'{-25'd68319}}, '{'{25'd669522}}, '{'{-25'd1544001}}, '{'{25'd1079434}}, '{'{25'd81982}}, '{'{-25'd1229735}}, '{'{-25'd109310}}, '{'{25'd232283}}, '{'{25'd628531}}, '{'{-25'd519221}}, '{'{-25'd341593}}, '{'{25'd1393700}}, '{'{-25'd1298054}}, '{'{25'd1448355}}, '{'{25'd1024779}}, '{'{-25'd1748957}}, '{'{-25'd655859}}, '{'{25'd1257062}}, '{'{-25'd1557664}}, '{'{-25'd478230}}, '{'{-25'd505558}}, '{'{25'd915469}}, '{'{25'd1544001}}, '{'{-25'd450903}}, '{'{25'd1298054}}},
    '{'{'{-25'd635322}}, '{'{-25'd698855}}, '{'{25'd1524774}}, '{'{-25'd1270645}}, '{'{25'd825919}}, '{'{25'd127064}}, '{'{-25'd762387}}, '{'{25'd762387}}, '{'{25'd698855}}, '{'{-25'd1016516}}, '{'{-25'd1143580}}, '{'{-25'd762387}}, '{'{25'd635322}}, '{'{25'd444726}}, '{'{25'd1334177}}, '{'{25'd1334177}}, '{'{-25'd952984}}, '{'{25'd1016516}}, '{'{25'd889451}}, '{'{25'd952984}}, '{'{25'd8068595}}, '{'{25'd571790}}, '{'{25'd1080048}}, '{'{-25'd635322}}, '{'{25'd1080048}}, '{'{-25'd127064}}, '{'{-25'd317661}}, '{'{25'd444726}}, '{'{25'd381193}}, '{'{-25'd1143580}}, '{'{-25'd1080048}}, '{'{-25'd1080048}}, '{'{-25'd1016516}}, '{'{25'd952984}}, '{'{-25'd127064}}, '{'{-25'd1016516}}, '{'{-25'd1207113}}, '{'{25'd952984}}, '{'{-25'd1016516}}, '{'{-25'd762387}}, '{'{-25'd1080048}}, '{'{-25'd127064}}, '{'{-25'd381193}}, '{'{25'd1016516}}, '{'{-25'd1397709}}, '{'{-25'd444726}}, '{'{-25'd317661}}, '{'{25'd762387}}, '{'{-25'd1461242}}, '{'{25'd889451}}, '{'{25'd571790}}, '{'{-25'd1270645}}, '{'{25'd889451}}, '{'{25'd1715371}}, '{'{-25'd698855}}, '{'{25'd1651838}}, '{'{-25'd889451}}, '{'{-25'd508258}}, '{'{-25'd1461242}}, '{'{25'd63532}}, '{'{-25'd1461242}}, '{'{-25'd2350693}}, '{'{25'd1715371}}, '{'{25'd1143580}}},
    '{'{'{-25'd925234}}, '{'{-25'd1206828}}, '{'{25'd295002}}, '{'{25'd335230}}, '{'{-25'd1367738}}, '{'{-25'd831370}}, '{'{25'd1381147}}, '{'{-25'd107274}}, '{'{-25'd1220237}}, '{'{25'd295002}}, '{'{-25'd1595694}}, '{'{25'd1622513}}, '{'{25'd362048}}, '{'{25'd1247055}}, '{'{-25'd1716377}}, '{'{-25'd1595694}}, '{'{25'd201138}}, '{'{-25'd107274}}, '{'{25'd67046}}, '{'{-25'd469322}}, '{'{25'd724097}}, '{'{-25'd402276}}, '{'{25'd1126372}}, '{'{-25'd563186}}, '{'{25'd1676149}}, '{'{25'd1314101}}, '{'{25'd1354329}}, '{'{-25'd750915}}, '{'{25'd160910}}, '{'{-25'd563186}}, '{'{25'd1542057}}, '{'{25'd1019099}}, '{'{25'd817961}}, '{'{-25'd348639}}, '{'{-25'd1582285}}, '{'{-25'd1582285}}, '{'{-25'd40228}}, '{'{-25'd1461602}}, '{'{-25'd791143}}, '{'{-25'd53637}}, '{'{25'd1072736}}, '{'{25'd1220237}}, '{'{-25'd898416}}, '{'{25'd992280}}, '{'{25'd1180009}}, '{'{-25'd1233646}}, '{'{-25'd67046}}, '{'{25'd348639}}, '{'{-25'd67046}}, '{'{-25'd1273874}}, '{'{-25'd683869}}, '{'{25'd630232}}, '{'{-25'd201138}}, '{'{-25'd831370}}, '{'{-25'd1193418}}, '{'{-25'd308411}}, '{'{25'd549777}}, '{'{25'd1542057}}, '{'{25'd281593}}, '{'{25'd737506}}, '{'{-25'd817961}}, '{'{25'd978871}}, '{'{-25'd1635922}}, '{'{25'd791143}}},
    '{'{'{25'd396779}}, '{'{25'd963605}}, '{'{-25'd207836}}, '{'{25'd2172836}}, '{'{25'd529038}}, '{'{-25'd1114759}}, '{'{25'd1587115}}, '{'{25'd566827}}, '{'{25'd623509}}, '{'{25'd774663}}, '{'{-25'd812452}}, '{'{25'd1719374}}, '{'{25'd755769}}, '{'{25'd793557}}, '{'{25'd566827}}, '{'{25'd226731}}, '{'{-25'd226731}}, '{'{-25'd1247019}}, '{'{-25'd1398173}}, '{'{-25'd566827}}, '{'{-25'd2418461}}, '{'{25'd1228125}}, '{'{25'd264519}}, '{'{-25'd831346}}, '{'{-25'd472356}}, '{'{-25'd1247019}}, '{'{25'd264519}}, '{'{25'd1001394}}, '{'{-25'd1039182}}, '{'{25'd1303701}}, '{'{25'd170048}}, '{'{25'd321202}}, '{'{25'd585721}}, '{'{25'd1662692}}, '{'{-25'd377884}}, '{'{25'd755769}}, '{'{25'd491250}}, '{'{25'd547933}}, '{'{25'd321202}}, '{'{25'd1662692}}, '{'{25'd94471}}, '{'{-25'd94471}}, '{'{25'd774663}}, '{'{-25'd1417067}}, '{'{25'd1624903}}, '{'{-25'd1133653}}, '{'{-25'd510144}}, '{'{25'd850240}}, '{'{-25'd434567}}, '{'{-25'd1549326}}, '{'{-25'd510144}}, '{'{-25'd56683}}, '{'{-25'd377884}}, '{'{-25'd1643798}}, '{'{25'd472356}}, '{'{25'd1360384}}, '{'{25'd1549326}}, '{'{-25'd188942}}, '{'{25'd1152548}}, '{'{25'd1001394}}, '{'{-25'd75577}}, '{'{-25'd113365}}, '{'{25'd944711}}, '{'{-25'd1322596}}},
    '{'{'{-25'd896018}}, '{'{25'd746682}}, '{'{25'd1393806}}, '{'{25'd1891594}}, '{'{25'd896018}}, '{'{25'd1294249}}, '{'{-25'd846240}}, '{'{25'd1443585}}, '{'{25'd1443585}}, '{'{-25'd1244470}}, '{'{-25'd1692479}}, '{'{-25'd1642700}}, '{'{25'd199115}}, '{'{-25'd199115}}, '{'{25'd348452}}, '{'{25'd149336}}, '{'{25'd1642700}}, '{'{-25'd597346}}, '{'{25'd348452}}, '{'{25'd2389382}}, '{'{-25'd6222350}}, '{'{25'd1443585}}, '{'{25'd1792037}}, '{'{25'd149336}}, '{'{25'd696903}}, '{'{-25'd448009}}, '{'{-25'd298673}}, '{'{-25'd647124}}, '{'{-25'd1194691}}, '{'{25'd6321908}}, '{'{-25'd2040931}}, '{'{25'd945797}}, '{'{25'd2140488}}, '{'{25'd1443585}}, '{'{25'd398230}}, '{'{-25'd149336}}, '{'{25'd199115}}, '{'{-25'd896018}}, '{'{-25'd49779}}, '{'{25'd1543143}}, '{'{-25'd597346}}, '{'{-25'd1045355}}, '{'{25'd696903}}, '{'{-25'd1642700}}, '{'{-25'd945797}}, '{'{-25'd1742258}}, '{'{-25'd547567}}, '{'{-25'd696903}}, '{'{-25'd1543143}}, '{'{25'd1244470}}, '{'{25'd796461}}, '{'{25'd2837392}}, '{'{25'd1144912}}, '{'{25'd448009}}, '{'{25'd2339604}}, '{'{-25'd398230}}, '{'{25'd597346}}, '{'{-25'd1443585}}, '{'{25'd995576}}, '{'{25'd945797}}, '{'{-25'd298673}}, '{'{-25'd746682}}, '{'{-25'd1294249}}, '{'{-25'd597346}}},
    '{'{'{25'd43650}}, '{'{-25'd873000}}, '{'{-25'd1615050}}, '{'{25'd698400}}, '{'{-25'd698400}}, '{'{-25'd1178550}}, '{'{25'd3535650}}, '{'{25'd785700}}, '{'{-25'd523800}}, '{'{25'd1353150}}, '{'{-25'd1658700}}, '{'{25'd305550}}, '{'{25'd654750}}, '{'{-25'd1615050}}, '{'{25'd785700}}, '{'{25'd1702350}}, '{'{25'd0}}, '{'{-25'd261900}}, '{'{25'd349200}}, '{'{25'd261900}}, '{'{-25'd2880900}}, '{'{25'd1396800}}, '{'{25'd2226150}}, '{'{-25'd1178550}}, '{'{-25'd1746000}}, '{'{-25'd218250}}, '{'{25'd1876950}}, '{'{25'd742050}}, '{'{-25'd523800}}, '{'{25'd2968200}}, '{'{-25'd567450}}, '{'{25'd261900}}, '{'{25'd2575350}}, '{'{-25'd392850}}, '{'{-25'd1091250}}, '{'{25'd1003950}}, '{'{-25'd2095200}}, '{'{25'd785700}}, '{'{-25'd305550}}, '{'{25'd742050}}, '{'{-25'd4845149}}, '{'{25'd611100}}, '{'{25'd261900}}, '{'{-25'd87300}}, '{'{25'd480150}}, '{'{-25'd130950}}, '{'{25'd829350}}, '{'{25'd829350}}, '{'{-25'd1396800}}, '{'{25'd829350}}, '{'{25'd742050}}, '{'{-25'd5587199}}, '{'{25'd218250}}, '{'{-25'd523800}}, '{'{25'd1091250}}, '{'{-25'd1134900}}, '{'{-25'd1222200}}, '{'{-25'd436500}}, '{'{25'd305550}}, '{'{25'd1353150}}, '{'{-25'd829350}}, '{'{25'd1964250}}, '{'{25'd130950}}, '{'{25'd1134900}}}
};
