localparam bit signed [0:2][0:26][19:0] Input0 = '{
    '{20'd44, -20'd81, -20'd11, 20'd64, -20'd61, 20'd123, 20'd67, -20'd25, -20'd119, 20'd83, -20'd107, 20'd114, -20'd92, -20'd41, -20'd58, 20'd88, -20'd40, 20'd12, -20'd70, 20'd65, 20'd102, -20'd89, -20'd41, 20'd46, -20'd40, -20'd47, 20'd37},
    '{-20'd103, -20'd51, -20'd56, -20'd119, 20'd20, -20'd13, 20'd80, 20'd115, 20'd69, 20'd126, -20'd49, 20'd47, 20'd64, -20'd46, -20'd29, 20'd88, 20'd49, 20'd115, -20'd99, 20'd19, 20'd19, 20'd14, 20'd39, -20'd96, 20'd65, -20'd119, 20'd57},
    '{-20'd1, -20'd96, -20'd97, 20'd74, 20'd116, 20'd23, 20'd35, 20'd126, 20'd75, -20'd14, 20'd55, -20'd100, -20'd94, 20'd0, 20'd0, 20'd36, -20'd75, 20'd5, -20'd90, 20'd104, 20'd116, -20'd111, -20'd49, 20'd4, -20'd23, -20'd86, 20'd58}
};
