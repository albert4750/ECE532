localparam bit signed [0:7][0:2][0:2][0:2][24:0] Weight1 = '{
    '{'{'{25'd1541, -25'd1228, -25'd2412}, '{25'd1251, 25'd893, 25'd1362}, '{25'd916, -25'd1139, 25'd2300}}, '{'{25'd826, 25'd2702, 25'd625}, '{25'd2836, 25'd2680, 25'd2657}, '{25'd2523, -25'd1876, -25'd1787}}, '{'{25'd2345, 25'd2233, -25'd514}, '{-25'd2256, -25'd1228, -25'd1251}, '{-25'd2323, 25'd1452, -25'd692}}},
    '{'{'{-25'd2286, 25'd1656, -25'd1557}, '{25'd1873, -25'd2346, 25'd2267}, '{25'd1695, -25'd2484, -25'd158}}, '{'{25'd848, -25'd867, -25'd256}, '{25'd631, 25'd1005, 25'd1301}, '{25'd1991, -25'd1557, -25'd2523}}, '{'{-25'd1577, -25'd2346, -25'd591}, '{-25'd848, -25'd1892, -25'd710}, '{-25'd1794, -25'd493, -25'd926}}},
    '{'{'{-25'd2705, 25'd195, 25'd307}, '{-25'd3290, 25'd3541, -25'd2398}, '{-25'd2844, 25'd362, -25'd1952}}, '{'{25'd1143, -25'd28, -25'd530}, '{25'd2008, 25'd3067, 25'd530}, '{25'd2649, 25'd976, -25'd1060}}, '{'{25'd1283, -25'd669, -25'd3234}, '{25'd3374, 25'd3541, 25'd2677}, '{25'd2398, 25'd3374, 25'd1645}}},
    '{'{'{25'd2496, -25'd930, 25'd1294}, '{25'd2701, 25'd1044, 25'd590}, '{25'd2882, 25'd1407, -25'd1861}}, '{'{25'd522, 25'd1770, 25'd1021}, '{-25'd2088, 25'd1679, -25'd2020}, '{-25'd2315, 25'd1906, 25'd2791}}, '{'{-25'd1225, 25'd1861, 25'd1906}, '{-25'd2156, -25'd658, -25'd1203}, '{25'd386, 25'd159, -25'd386}}},
    '{'{'{25'd1663, -25'd1422, -25'd963}, '{-25'd2778, -25'd700, 25'd2100}, '{25'd963, 25'd1510, -25'd2669}}, '{'{25'd22, -25'd109, 25'd1006}, '{-25'd2603, 25'd1860, -25'd1685}, '{25'd131, -25'd2560, -25'd2078}}, '{'{-25'd809, 25'd2560, 25'd1378}, '{25'd0, -25'd2210, -25'd350}, '{25'd853, 25'd2035, -25'd634}}},
    '{'{'{-25'd1373, -25'd824, -25'd23}, '{-25'd984, 25'd503, 25'd1968}, '{25'd503, -25'd458, 25'd1464}}, '{'{25'd46, 25'd1487, -25'd2563}, '{-25'd1190, 25'd69, -25'd1281}, '{25'd1922, 25'd1739, 25'd1281}}, '{'{-25'd686, -25'd1991, -25'd1808}, '{25'd1968, 25'd2906, 25'd1167}, '{25'd1281, 25'd847, 25'd2082}}},
    '{'{'{25'd1762, -25'd655, 25'd1920}, '{25'd632, 25'd1175, 25'd2259}, '{25'd1288, 25'd1581, 25'd2123}}, '{'{-25'd1265, 25'd904, -25'd2891}, '{25'd2056, -25'd2372, 25'd1175}, '{-25'd2078, -25'd1536, 25'd203}}, '{'{25'd1807, -25'd2440, 25'd994}, '{-25'd2869, -25'd1152, -25'd1084}, '{-25'd2236, -25'd181, -25'd2214}}},
    '{'{'{25'd870, 25'd2154, -25'd653}, '{25'd1610, -25'd1284, 25'd2219}, '{-25'd435, -25'd196, 25'd1784}}, '{'{25'd1762, -25'd500, -25'd239}, '{-25'd413, 25'd653, -25'd1371}, '{-25'd1871, 25'd1719, -25'd2437}}, '{'{-25'd370, 25'd2763, -25'd805}, '{25'd2524, 25'd1066, 25'd1436}, '{25'd935, 25'd2197, -25'd914}}}
};
