localparam bit signed [0:10][15:0] Output7 = '{16'd8616, -16'd24872, 16'd12842, -16'd4887, 16'd18550, 16'd21168, 16'd17341, -16'd15137, 16'd1429, -16'd27696, -16'd12814};
