localparam bit signed [0:15][7:0] Output7 = '{38, 75, -9, -4, -84, 69, -2, -96, -90, 31, -66, -97, -95, -88, -63, -79};
