localparam bit signed [0:7][35:0] Bias2 = '{36'd0, 36'd0, 36'd0, 36'd0, 36'd0, 36'd0, 36'd0, 36'd0};
