localparam bit signed [0:10][36:0] Bias = '{-37'd12125, -37'd20934, -37'd15439, 37'd29802, -37'd24375, 37'd23852, -37'd14579, 37'd15225, -37'd30906, 37'd8742, 37'd3751};
