localparam bit signed [0:15][7:0] Output1 = '{-54, -122, -28, -24, -48, -14, 17, 13, -89, -48, -74, -38, 68, 98, -101, 57};
