localparam bit signed [0:26][19:0] Output7 = '{-20'd156, 20'd125, 20'd71, -20'd98, 20'd2, 20'd145, -20'd66, 20'd123, -20'd262, -20'd50, -20'd44, 20'd11, 20'd15, 20'd76, -20'd289, 20'd150, -20'd8, 20'd104, 20'd115, -20'd23, -20'd40, -20'd295, -20'd119, -20'd44, 20'd155, -20'd30, 20'd2};
