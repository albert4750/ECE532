localparam bit signed [0:7][0:2][0:2][0:2][19:0] Weight1 = '{
    '{'{'{20'd38994, -20'd50795, 20'd37455}, '{20'd8209, 20'd30785, 20'd26680}, '{20'd65161, -20'd18984, 20'd1539}}, '{'{20'd14366, 20'd49769, 20'd10262}, '{-20'd7696, -20'd48743, -20'd7696}, '{-20'd9235, -20'd8722, -20'd23602}}, '{'{20'd51821, 20'd31298, -20'd26680}, '{20'd34889, -20'd15905, -20'd18984}, '{20'd3592, 20'd0, 20'd22062}}},
    '{'{'{20'd14526, -20'd9338, -20'd66405}, '{20'd0, -20'd39947, 20'd58623}, '{20'd42022, 20'd14526, -20'd22827}}, '{'{20'd2594, -20'd10376, 20'd24902}, '{-20'd18676, -20'd33721, -20'd20751}, '{-20'd7263, 20'd35796, -20'd26458}}, '{'{20'd2075, -20'd25421, -20'd47210}, '{-20'd42022, -20'd519, -20'd20233}, '{-20'd17639, -20'd28015, 20'd6225}}},
    '{'{'{20'd42128, 20'd53868, -20'd33840}, '{20'd8287, 20'd51796, -20'd691}, '{20'd26934, -20'd28315, -20'd15194}}, '{'{20'd56631, -20'd66990, 20'd22790}, '{20'd81493, 20'd85636, 20'd15194}, '{-20'd15194, 20'd55940, -20'd2762}}, '{'{20'd26243, 20'd15194, -20'd35221}, '{20'd44890, -20'd21409, -20'd7597}, '{-20'd62155, -20'd87708, -20'd14503}}},
    '{'{'{-20'd9827, -20'd8793, -20'd43963}, '{20'd32067, 20'd51204, 20'd56376}, '{-20'd66203, 20'd8275, -20'd61031}}, '{'{-20'd24309, 20'd13448, -20'd66203}, '{20'd48101, 20'd45515, -20'd5689}, '{-20'd47584, 20'd56376, -20'd65169}}, '{'{-20'd51204, 20'd17585, -20'd517}, '{20'd12930, 20'd56894, 20'd26895}, '{20'd18102, -20'd23275, -20'd32584}}},
    '{'{'{-20'd15069, -20'd18187, -20'd50923}, '{20'd36373, -20'd43129, -20'd520}, '{-20'd33256, -20'd11432, 20'd11432}}, '{'{20'd23903, -20'd48325, 20'd21304}, '{-20'd53001, -20'd22344, 20'd25981}, '{20'd19746, 20'd18187, -20'd66512}}, '{'{20'd22863, 20'd15589, 20'd18706}, '{-20'd29099, -20'd48844, -20'd56119}, '{-20'd44168, 20'd25981, 20'd19226}}},
    '{'{'{-20'd45195, -20'd36587, 20'd41967}, '{-20'd3228, 20'd45195, 20'd8609}, '{20'd7533, 20'd53804, 20'd8609}}, '{'{-20'd137739, -20'd3228, 20'd25826}, '{-20'd112989, -20'd2152, -20'd22598}, '{-20'd36587, 20'd45195, -20'd49500}}, '{'{-20'd54880, 20'd67793, -20'd50576}, '{-20'd99000, -20'd21522, -20'd54880}, '{-20'd22598, 20'd74250, 20'd3228}}},
    '{'{'{20'd14295, 20'd25731, -20'd33355}, '{20'd68616, 20'd78146, 20'd74334}, '{20'd121031, 20'd38120, -20'd20013}}, '{'{20'd36214, -20'd17154, -20'd8577}, '{-20'd1906, 20'd61945, 20'd66710}, '{-20'd40026, 20'd51462, -20'd45744}}, '{'{20'd65757, 20'd0, -20'd17154}, '{-20'd7624, 20'd13342, -20'd40979}, '{-20'd25731, 20'd49556, -20'd28590}}},
    '{'{'{20'd6436, 20'd2861, -20'd47201}, '{20'd38619, -20'd25746, 20'd13588}, '{-20'd17164, -20'd21455, -20'd25746}}, '{'{20'd8582, 20'd67940, 20'd24316}, '{20'd76522, 20'd27891, -20'd7867}, '{20'd38619, 20'd43625, 20'd33613}}, '{'{-20'd36473, 20'd13588, -20'd36473}, '{-20'd2861, 20'd90826, 20'd65795}, '{20'd22170, 20'd55783, -20'd21455}}}
};
