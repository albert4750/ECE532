logic signed [7:0] convolve23_weight[4][8][3][3] = '{
    '{
        '{'{-113, 101, 105}, '{-11, 92, -37}, '{55, 59, 123}},
        '{'{109, 55, -3}, '{33, -117, -1}, '{91, -94, 88}},
        '{'{-115, 7, 24}, '{65, -29, -46}, '{-18, -88, 55}},
        '{'{-63, 106, -101}, '{15, 15, -87}, '{77, -122, -2}},
        '{'{122, 96, 92}, '{-72, 52, 6}, '{-50, 31, 6}},
        '{'{-95, -1, 58}, '{122, -2, -82}, '{-1, -102, -77}},
        '{'{32, 60, 123}, '{-82, -33, 7}, '{49, -89, 65}},
        '{'{-123, -27, 27}, '{38, -83, 23}, '{-116, 9, 29}}
    },
    '{
        '{'{29, -115, -41}, '{-104, 9, -60}, '{37, 56, 75}},
        '{'{-42, 60, 24}, '{-27, -24, 104}, '{52, -75, -30}},
        '{'{46, 33, 122}, '{13, 97, 71}, '{-116, 73, 46}},
        '{'{-99, -116, 55}, '{-80, 118, -93}, '{-94, -70, 60}},
        '{'{1, 17, 43}, '{112, 55, -119}, '{55, 121, 125}},
        '{'{16, -61, 41}, '{86, -81, 84}, '{-40, 97, 123}},
        '{'{-70, 84, 85}, '{-92, 108, -116}, '{-102, -126, 122}},
        '{'{122, -106, -82}, '{-45, 121, -110}, '{-94, -33, 67}}
    },
    '{
        '{'{-128, 27, -80}, '{110, 86, 116}, '{3, 124, 96}},
        '{'{-117, -16, 88}, '{28, -88, 73}, '{-126, 78, -69}},
        '{'{116, -118, 4}, '{73, -19, -1}, '{-38, -21, 125}},
        '{'{-120, -91, 104}, '{98, 108, 118}, '{-26, -37, 112}},
        '{'{58, 58, 49}, '{117, -109, -93}, '{36, -4, -54}},
        '{'{-79, 18, -124}, '{88, 79, -79}, '{94, -115, 51}},
        '{'{16, 55, -24}, '{109, 75, -67}, '{-30, -111, 70}},
        '{'{-104, -35, 93}, '{-62, 75, 122}, '{-82, 40, 81}}
    },
    '{
        '{'{39, 127, -119}, '{-21, -102, -108}, '{57, 68, -22}},
        '{'{-62, -76, -89}, '{-45, 63, -12}, '{7, -97, -32}},
        '{'{68, 116, 27}, '{24, 106, -73}, '{8, -84, -75}},
        '{'{90, -90, 27}, '{98, -85, 76}, '{111, -120, 40}},
        '{'{-8, 109, -96}, '{64, 111, 81}, '{76, -112, -11}},
        '{'{120, -53, -49}, '{92, -77, 64}, '{-18, 92, 36}},
        '{'{-68, -110, 81}, '{25, -88, 25}, '{-124, 10, -31}},
        '{'{-42, 97, -18}, '{82, 35, 112}, '{-44, 5, -70}}
    }
};
