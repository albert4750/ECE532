wire signed [7:0] convolve0_weight[4][3][3][3];
assign convolve0_weight = '{'{'{'{44, -81, -11}, '{64, -61, 123}, '{67, -25, -119}}, '{'{83, -107, 114}, '{-92, -41, -58}, '{88, -40, 12}}, '{'{-70, 65, 102}, '{-89, -41, 46}, '{-40, -47, 37}}}, '{'{'{-103, -51, -56}, '{-119, 20, -13}, '{80, 115, 69}}, '{'{126, -49, 47}, '{64, -46, -29}, '{88, 49, 115}}, '{'{-99, 19, 19}, '{14, 39, -96}, '{65, -119, 57}}}, '{'{'{-1, -96, -97}, '{74, 116, 23}, '{35, 126, 75}}, '{'{-14, 55, -100}, '{-94, 0, 0}, '{36, -75, 5}}, '{'{-90, 104, 116}, '{-111, -49, 4}, '{-23, -86, 58}}}, '{'{'{-97, -8, -127}, '{-63, 103, 41}, '{-71, -93, -26}}, '{'{-9, -117, 46}, '{-46, -37, 0}, '{14, -29, -75}}, '{'{12, -7, 42}, '{-44, 75, -60}, '{-122, 68, -81}}}};
