localparam bit signed [0:7][47:0] Bias1 = '{-48'd33184, -48'd572822, 48'd299697, -48'd44335, -48'd408385, 48'd116897, -48'd14847, -48'd110936};
