localparam bit signed [0:2][0:26][19:0] Input6 = '{
    '{-20'd76, 20'd110, 20'd49, 20'd91, -20'd77, 20'd99, -20'd23, -20'd110, -20'd11, -20'd94, -20'd77, 20'd30, 20'd53, -20'd70, 20'd43, -20'd73, 20'd124, 20'd124, -20'd110, 20'd45, -20'd41, 20'd65, -20'd58, 20'd106, -20'd75, -20'd80, -20'd34},
    '{-20'd69, -20'd48, 20'd26, -20'd4, 20'd35, -20'd70, 20'd49, -20'd22, 20'd73, -20'd84, -20'd115, -20'd7, -20'd58, -20'd90, 20'd39, 20'd8, -20'd115, 20'd120, 20'd7, 20'd80, 20'd120, -20'd106, 20'd120, -20'd49, 20'd89, -20'd120, 20'd99},
    '{-20'd122, 20'd81, 20'd71, 20'd84, 20'd89, 20'd66, -20'd68, 20'd16, -20'd72, -20'd14, 20'd109, 20'd23, -20'd104, -20'd124, -20'd28, 20'd108, -20'd79, -20'd41, -20'd98, -20'd74, 20'd25, -20'd108, -20'd31, -20'd27, 20'd57, 20'd23, 20'd27}
};
