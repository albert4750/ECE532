localparam bit signed [0:2][47:0] Bias3 = '{48'd228235, -48'd340770, 48'd770915};
