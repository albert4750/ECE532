localparam bit signed [0:10][15:0] Output9 = '{16'd2749, 16'd12041, 16'd24487, 16'd14562, -16'd19280, -16'd713, 16'd20377, -16'd8372, 16'd25238, 16'd28073, -16'd11913};
