localparam bit signed [0:31][47:0] Bias2 = '{-48'd52399, -48'd155244, -48'd130475, 48'd35991, 48'd145531, 48'd37959, -48'd108128, 48'd12086, 48'd28740, 48'd38917, 48'd41685, -48'd69134, 48'd114614, -48'd103098, 48'd161566, 48'd75549, 48'd126360, 48'd144386, -48'd42682, 48'd2957, -48'd3901, -48'd18621, 48'd37921, 48'd126545, -48'd148717, 48'd149139, 48'd155937, -48'd45224, 48'd89389, 48'd42271, -48'd66330, -48'd137843};
