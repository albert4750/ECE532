localparam bit signed [0:31][47:0] Bias2 = '{48'd2836, 48'd2744, 48'd2376, 48'd2517, 48'd2806, 48'd2262, 48'd3102, -48'd4180, 48'd3053, 48'd3013, 48'd3213, 48'd3616, 48'd3526, 48'd3128, 48'd3399, 48'd2162, 48'd1801, 48'd2248, -48'd1873, 48'd2868, 48'd3621, 48'd2809, 48'd1078, 48'd2444, 48'd2699, 48'd3371, 48'd3883, 48'd1535, 48'd2348, 48'd2224, 48'd2403, 48'd3596};
