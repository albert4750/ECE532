localparam bit signed [0:46][15:0] Input3 = '{-16'd30464, -16'd20859, 16'd3419, 16'd1131, -16'd1122, -16'd18487, -16'd14381, 16'd28167, 16'd27797, 16'd10213, -16'd8740, -16'd19064, 16'd18091, -16'd22994, -16'd24576, -16'd25240, 16'd691, 16'd13862, 16'd29785, -16'd5046, -16'd13837, -16'd5406, -16'd30085, -16'd7849, -16'd17312, -16'd25773, -16'd3814, 16'd23246, -16'd26592, -16'd5005, 16'd6598, -16'd26783, 16'd4524, 16'd827, -16'd22727, 16'd23218, -16'd22355, -16'd2327, -16'd29564, 16'd28089, -16'd32675, 16'd15707, -16'd19055, 16'd2467, 16'd3778, -16'd32364, -16'd27731};
