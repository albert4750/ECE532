localparam bit signed [0:63][0:2][0:8][0:8][24:0] Weight1 = '{
    '{'{'{25'd9604, 25'd3078, 25'd11327, -25'd5417, 25'd13297, 25'd8865, 25'd3078, 25'd13543, 25'd12558}, '{25'd5048, 25'd4432, -25'd2955, -25'd3201, -25'd8988, -25'd862, -25'd1847, -25'd7387, 25'd8249}, '{25'd11820, -25'd8742, -25'd7757, 25'd9480, 25'd7757, 25'd13174, 25'd13667, -25'd6156, 25'd9111}, '{25'd2462, -25'd3694, 25'd13543, 25'd0, 25'd9850, 25'd1477, -25'd7757, 25'd6649, 25'd12189}, '{-25'd5664, -25'd4309, 25'd9973, -25'd9604, 25'd2093, 25'd246, 25'd4063, 25'd15637, 25'd1970}, '{25'd5294, 25'd4925, 25'd3694, -25'd9111, 25'd1970, 25'd6279, 25'd5787, 25'd9727, 25'd1477}, '{-25'd616, 25'd9111, -25'd492, -25'd5417, 25'd13913, -25'd5048, 25'd616, 25'd12435, 25'd862}, '{25'd10342, -25'd3078, 25'd8742, -25'd1724, 25'd1354, 25'd13174, -25'd5540, -25'd1108, 25'd6649}, '{-25'd4186, -25'd1231, -25'd1970, 25'd4432, 25'd6033, 25'd11943, 25'd6649, 25'd13790, 25'd15144}}, '{'{25'd985, -25'd2832, 25'd1354, -25'd1970, -25'd7264, -25'd12189, -25'd862, -25'd3324, 25'd3201}, '{-25'd11573, -25'd8495, -25'd246, -25'd2709, 25'd9604, 25'd5540, 25'd9234, -25'd11327, -25'd8988}, '{-25'd12312, -25'd11573, -25'd2093, -25'd1354, -25'd3571, 25'd8126, 25'd369, -25'd5540, 25'd6525}, '{25'd6402, 25'd5910, 25'd4925, -25'd1601, 25'd8988, 25'd5048, 25'd6402, -25'd3940, -25'd12805}, '{25'd6649, -25'd11204, -25'd10096, -25'd12189, -25'd8742, -25'd11204, -25'd6895, -25'd3694, -25'd11081}, '{-25'd10589, -25'd2709, 25'd7757, -25'd5787, -25'd8619, -25'd10342, 25'd8249, -25'd12805, -25'd3201}, '{-25'd2955, 25'd3940, -25'd5540, -25'd8495, -25'd9604, -25'd3447, -25'd7141, -25'd6402, -25'd9604}, '{25'd8003, -25'd11327, -25'd2955, -25'd10835, -25'd2216, -25'd492, 25'd3447, -25'd9850, -25'd11697}, '{-25'd4186, -25'd3078, -25'd11820, 25'd9727, 25'd8988, -25'd5417, 25'd5910, -25'd6402, -25'd4556}}, '{'{-25'd7018, 25'd5417, -25'd9604, -25'd2462, 25'd4309, -25'd4802, 25'd2832, -25'd10096, -25'd8619}, '{-25'd10835, 25'd2216, -25'd7510, -25'd3817, -25'd9480, 25'd10096, 25'd9850, -25'd8249, -25'd2093}, '{-25'd616, -25'd7880, -25'd2709, -25'd5910, 25'd9973, 25'd1108, -25'd4556, 25'd862, 25'd1231}, '{-25'd2709, 25'd11697, 25'd1231, 25'd739, 25'd8003, -25'd1231, 25'd9604, -25'd4432, 25'd2216}, '{25'd6649, 25'd6156, 25'd9604, -25'd6649, 25'd8865, -25'd10096, -25'd3817, 25'd1108, -25'd2586}, '{-25'd6033, -25'd246, -25'd10096, -25'd4309, 25'd369, -25'd10835, 25'd8249, -25'd5540, -25'd1847}, '{-25'd9727, -25'd739, -25'd10835, -25'd6156, 25'd5787, -25'd10589, 25'd2586, 25'd10096, 25'd11204}, '{-25'd1108, -25'd8495, 25'd2955, 25'd8495, -25'd1970, 25'd246, 25'd369, -25'd1354, -25'd369}, '{25'd12312, -25'd1970, -25'd5294, 25'd10958, -25'd11327, 25'd12189, 25'd4679, -25'd3078, 25'd4802}}},
    '{'{'{25'd0, 25'd6256, 25'd7277, -25'd12257, 25'd2426, -25'd9831, 25'd3064, 25'd10469, 25'd10725}, '{25'd2681, -25'd3703, -25'd6639, -25'd3064, -25'd2554, 25'd10980, 25'd9320, -25'd3447, -25'd3192}, '{-25'd12512, -25'd13278, 25'd2554, 25'd8427, -25'd5107, 25'd3958, -25'd4086, -25'd4341, 25'd9065}, '{25'd1149, 25'd6001, -25'd1532, 25'd1277, 25'd7533, -25'd13278, -25'd3703, 25'd3703, 25'd2681}, '{-25'd11363, -25'd10597, -25'd9448, -25'd8171, -25'd3575, -25'd12895, -25'd2170, 25'd8937, 25'd5235}, '{25'd9448, -25'd10469, -25'd7277, -25'd9193, -25'd7661, -25'd1660, 25'd3064, 25'd638, 25'd8937}, '{-25'd4724, -25'd5618, 25'd128, -25'd7916, -25'd16215, -25'd3064, -25'd7661, -25'd4852, -25'd8171}, '{25'd6639, -25'd7277, -25'd13534, -25'd6256, -25'd10597, -25'd14683, 25'd8299, -25'd8299, 25'd8044}, '{-25'd5107, -25'd8427, -25'd4979, -25'd9576, 25'd5107, 25'd383, -25'd11491, 25'd11108, 25'd2554}}, '{'{25'd8427, 25'd8427, 25'd6767, -25'd8299, 25'd1915, 25'd2937, -25'd766, -25'd1660, 25'd1660}, '{-25'd8427, 25'd8044, 25'd1915, -25'd8044, -25'd9703, -25'd5745, -25'd8682, 25'd8937, 25'd5107}, '{25'd4086, 25'd12257, 25'd1404, 25'd4341, -25'd7661, -25'd128, -25'd6639, 25'd10597, 25'd9065}, '{25'd4852, 25'd894, 25'd8171, 25'd11746, 25'd8937, 25'd8810, 25'd8937, -25'd9320, 25'd7150}, '{-25'd4086, 25'd6511, -25'd9320, 25'd11618, 25'd12768, 25'd383, -25'd7150, -25'd7277, 25'd1915}, '{-25'd766, 25'd4852, 25'd6767, -25'd7533, 25'd128, -25'd8299, -25'd8299, -25'd7533, -25'd8299}, '{-25'd6256, -25'd7022, -25'd7277, 25'd3575, 25'd4596, -25'd1277, 25'd7022, 25'd766, -25'd766}, '{-25'd3192, 25'd10469, 25'd7661, 25'd11235, -25'd7150, -25'd638, 25'd12640, 25'd128, -25'd4341}, '{25'd7788, 25'd5873, -25'd2043, 25'd9065, 25'd12385, -25'd6256, -25'd9576, -25'd10214, -25'd7661}}, '{'{25'd1404, 25'd3320, 25'd5490, 25'd10214, 25'd10086, -25'd4469, 25'd8171, -25'd9065, 25'd7661}, '{25'd3703, 25'd9576, 25'd8299, 25'd11618, 25'd3575, 25'd1021, 25'd11618, 25'd255, -25'd3703}, '{25'd638, 25'd2043, 25'd9065, -25'd10342, -25'd3447, 25'd11874, 25'd5362, 25'd4724, 25'd3447}, '{25'd0, -25'd1915, 25'd12512, 25'd6767, -25'd3192, 25'd10214, 25'd8937, 25'd5362, 25'd7022}, '{25'd3958, 25'd1532, 25'd9703, -25'd5490, -25'd4086, 25'd1660, 25'd1277, 25'd12129, 25'd3320}, '{25'd6256, -25'd8810, -25'd10214, 25'd9831, 25'd11235, -25'd10469, -25'd5745, 25'd5362, 25'd7533}, '{-25'd3575, 25'd8937, -25'd1915, 25'd4086, 25'd9959, 25'd9320, 25'd9320, -25'd8937, 25'd7533}, '{-25'd8937, 25'd9320, 25'd6639, -25'd7022, 25'd128, 25'd1660, 25'd6128, -25'd5235, 25'd8682}, '{-25'd10086, -25'd10469, 25'd9959, -25'd5490, -25'd1277, -25'd11363, -25'd7022, -25'd766, -25'd7916}}},
    '{'{'{25'd10553, -25'd5965, 25'd2294, -25'd6118, 25'd7953, -25'd4436, 25'd3365, -25'd9483, -25'd14224}, '{-25'd2294, -25'd6271, 25'd4588, 25'd10248, -25'd6577, 25'd11012, -25'd7647, -25'd1988, 25'd1529}, '{25'd11777, 25'd11777, 25'd9942, 25'd6271, 25'd11318, -25'd10248, 25'd6271, -25'd7953, 25'd7953}, '{-25'd765, 25'd7953, -25'd7953, -25'd6730, 25'd11624, -25'd6577, -25'd3365, -25'd11318, -25'd12389}, '{25'd7189, 25'd14377, -25'd6730, 25'd13918, -25'd7036, 25'd2447, 25'd153, 25'd2753, -25'd13001}, '{25'd1988, 25'd8259, -25'd612, 25'd11471, -25'd12083, -25'd4283, -25'd3518, -25'd14377, 25'd153}, '{25'd10248, 25'd6271, -25'd6271, -25'd3977, -25'd11777, -25'd13460, -25'd9636, -25'd19577, -25'd15601}, '{-25'd5506, 25'd7495, 25'd1682, -25'd12236, -25'd11777, -25'd3059, 25'd5506, -25'd9942, -25'd13460}, '{25'd6883, -25'd8718, 25'd153, -25'd6271, 25'd153, 25'd3977, 25'd6730, -25'd13154, -25'd13001}}, '{'{-25'd9330, -25'd4436, -25'd10248, 25'd459, 25'd1835, 25'd1682, 25'd2753, 25'd2753, 25'd4894}, '{25'd9330, -25'd2294, -25'd1071, 25'd5659, 25'd9942, -25'd10553, -25'd10706, 25'd4436, 25'd1377}, '{25'd6577, 25'd5047, 25'd3365, -25'd4588, 25'd7495, 25'd0, 25'd8871, 25'd6730, -25'd14989}, '{25'd9330, 25'd6271, 25'd5812, 25'd9636, 25'd8412, 25'd2753, -25'd3059, 25'd1529, -25'd1377}, '{-25'd7953, -25'd12695, 25'd5353, 25'd5965, -25'd612, 25'd3671, 25'd1377, 25'd3212, -25'd4130}, '{-25'd1224, -25'd5047, 25'd0, -25'd4894, 25'd4588, 25'd3365, -25'd10401, 25'd306, -25'd3518}, '{-25'd6883, 25'd8106, -25'd8871, 25'd2906, -25'd8412, 25'd7647, -25'd9483, -25'd10553, -25'd7342}, '{-25'd5506, -25'd11624, -25'd10095, -25'd11012, 25'd8259, 25'd3518, 25'd1377, -25'd14071, 25'd5965}, '{25'd3059, -25'd8718, 25'd4588, -25'd8871, -25'd11318, 25'd153, -25'd6730, 25'd7189, -25'd1988}}, '{'{25'd6424, 25'd1071, -25'd5659, -25'd7953, 25'd1377, 25'd12083, -25'd2294, 25'd2447, -25'd765}, '{25'd5353, 25'd3977, 25'd7495, 25'd6271, 25'd11777, -25'd7647, 25'd10553, 25'd2753, 25'd6424}, '{-25'd3518, 25'd11777, 25'd15142, -25'd7495, 25'd612, -25'd9024, 25'd6577, 25'd2600, 25'd2141}, '{25'd5353, -25'd5965, -25'd7495, 25'd4588, -25'd3365, 25'd4130, -25'd6424, 25'd9024, -25'd7953}, '{-25'd3671, 25'd10248, -25'd5353, 25'd1377, -25'd5353, 25'd10095, 25'd12695, -25'd2447, -25'd9483}, '{25'd11777, -25'd1071, 25'd11012, 25'd3212, 25'd4588, -25'd5506, -25'd7495, 25'd7953, 25'd13154}, '{-25'd1071, 25'd5812, -25'd7189, -25'd6118, -25'd306, -25'd3059, 25'd11624, 25'd7036, -25'd10401}, '{25'd11777, 25'd10248, -25'd8259, 25'd2447, -25'd1682, 25'd9636, 25'd8259, -25'd2447, -25'd918}, '{25'd6118, 25'd9024, 25'd6577, -25'd6424, 25'd9789, -25'd5047, -25'd1682, 25'd7036, 25'd11012}}},
    '{'{'{-25'd4138, -25'd2633, 25'd7523, -25'd8275, 25'd7523, 25'd7711, -25'd2633, 25'd13165, 25'd3573}, '{25'd13165, 25'd6018, 25'd1128, 25'd3950, -25'd8275, -25'd8275, -25'd7335, -25'd3950, -25'd9968}, '{-25'd10908, 25'd1505, 25'd6583, -25'd5266, -25'd12413, -25'd8651, -25'd10532, 25'd4702, 25'd752}, '{-25'd5266, 25'd1128, 25'd10156, -25'd12601, 25'd9028, 25'd9028, -25'd4890, -25'd9216, 25'd1128}, '{-25'd7899, -25'd4326, 25'd9216, -25'd10720, -25'd5454, 25'd6395, 25'd6959, 25'd564, -25'd7147}, '{25'd1317, -25'd12789, -25'd4514, 25'd2445, -25'd4514, -25'd9404, -25'd12789, 25'd10720, -25'd1128}, '{25'd9592, -25'd564, -25'd1505, 25'd376, 25'd2257, -25'd13165, -25'd3761, 25'd564, -25'd2445}, '{25'd7899, 25'd8087, -25'd564, -25'd14482, -25'd5454, 25'd8087, 25'd2257, -25'd11284, -25'd11849}, '{-25'd15986, -25'd12225, -25'd15046, -25'd5266, -25'd6018, -25'd4138, -25'd9780, -25'd8087, 25'd4514}}, '{'{25'd5266, -25'd376, -25'd4514, -25'd14670, 25'd4514, -25'd16551, 25'd3573, -25'd1693, 25'd4138}, '{-25'd11849, -25'd6959, -25'd6583, -25'd18807, -25'd16174, -25'd11284, -25'd16362, -25'd15610, -25'd15046}, '{-25'd14858, -25'd16551, -25'd17303, 25'd376, 25'd1881, -25'd4702, -25'd7335, -25'd7523, -25'd1505}, '{-25'd10532, 25'd2633, 25'd0, -25'd19184, -25'd10156, 25'd2633, -25'd11473, -25'd17115, -25'd15610}, '{-25'd5830, -25'd4326, -25'd12977, -25'd18807, -25'd13541, -25'd376, -25'd6771, -25'd11096, -25'd8275}, '{-25'd3009, 25'd188, -25'd18431, -25'd1505, -25'd18619, -25'd16551, -25'd18807, -25'd17115, -25'd5078}, '{-25'd1505, 25'd1128, -25'd21252, -25'd13729, -25'd9028, 25'd752, -25'd5266, -25'd1317, -25'd564}, '{-25'd3385, -25'd3197, -25'd6583, -25'd4702, -25'd4326, -25'd4138, -25'd9216, -25'd3009, -25'd9592}, '{-25'd4890, -25'd10908, -25'd15046, -25'd24074, -25'd21441, -25'd22381, -25'd9968, 25'd1317, -25'd5454}}, '{'{25'd12601, 25'd5454, -25'd5830, 25'd7147, 25'd940, -25'd376, 25'd11284, 25'd3573, 25'd3009}, '{25'd376, 25'd14294, 25'd9404, -25'd4702, -25'd7711, 25'd1317, 25'd9592, -25'd1505, -25'd6959}, '{25'd7711, 25'd7899, 25'd11661, 25'd6959, 25'd9780, 25'd10344, 25'd7523, 25'd9404, 25'd14294}, '{25'd10156, -25'd376, -25'd3950, -25'd2069, 25'd12037, -25'd7147, 25'd15986, -25'd4702, 25'd12977}, '{25'd2445, 25'd13353, 25'd9592, -25'd1317, -25'd3009, 25'd11284, 25'd9968, 25'd1317, -25'd7335}, '{25'd11849, 25'd3009, -25'd2069, -25'd7899, 25'd7523, 25'd11284, 25'd5078, 25'd4702, 25'd9968}, '{25'd5830, 25'd5830, 25'd5830, 25'd2821, 25'd12601, -25'd5078, 25'd9404, 25'd11661, -25'd7899}, '{-25'd6959, -25'd2257, 25'd6395, 25'd9968, 25'd4326, -25'd2257, -25'd5454, -25'd376, 25'd8840}, '{25'd4138, 25'd5454, -25'd10156, -25'd6018, 25'd7899, -25'd8651, 25'd4514, -25'd9592, -25'd10156}}},
    '{'{'{-25'd12734, -25'd4825, 25'd536, -25'd7372, 25'd2547, -25'd2145, 25'd10857, 25'd5630, 25'd6836}, '{25'd3083, -25'd4021, -25'd6702, 25'd3485, -25'd8042, 25'd2279, 25'd7104, -25'd5362, 25'd7238}, '{-25'd10455, -25'd11662, -25'd9651, -25'd12466, 25'd268, 25'd10723, -25'd7372, -25'd7908, 25'd3083}, '{25'd4289, -25'd3887, 25'd5630, -25'd402, -25'd4155, 25'd4021, -25'd3887, 25'd4960, 25'd4557}, '{-25'd10187, 25'd5630, -25'd12466, -25'd1206, -25'd7908, 25'd11393, 25'd2681, -25'd10187, -25'd9115}, '{-25'd11930, 25'd3753, -25'd9919, 25'd4289, -25'd1877, 25'd402, -25'd8311, -25'd5764, 25'd134}, '{-25'd4691, -25'd8713, -25'd5898, -25'd11125, 25'd4289, 25'd9919, 25'd2949, -25'd5362, -25'd1340}, '{25'd4557, -25'd2279, -25'd536, -25'd6300, 25'd9383, 25'd11796, 25'd8311, -25'd4960, 25'd12064}, '{-25'd11528, -25'd8311, 25'd1743, -25'd8713, -25'd268, 25'd2949, -25'd5094, -25'd8713, -25'd9249}}, '{'{-25'd4960, 25'd8042, -25'd2145, 25'd6702, -25'd9517, -25'd2413, 25'd2413, -25'd1474, -25'd8311}, '{-25'd2547, -25'd6166, -25'd6568, 25'd6300, -25'd10723, -25'd5630, 25'd3351, -25'd134, 25'd8311}, '{-25'd14074, -25'd804, 25'd8311, 25'd3485, -25'd2815, 25'd3083, 25'd4021, 25'd134, 25'd13940}, '{-25'd14074, -25'd12198, 25'd10455, 25'd5228, -25'd6032, 25'd9651, -25'd3217, 25'd10723, 25'd11796}, '{-25'd4557, -25'd2815, 25'd10589, -25'd11393, 25'd4155, -25'd8445, 25'd7104, -25'd1743, 25'd6032}, '{25'd6970, 25'd1474, -25'd1743, 25'd3619, -25'd9785, -25'd3753, -25'd3217, 25'd5496, 25'd4557}, '{-25'd9249, 25'd11528, 25'd8445, 25'd10589, 25'd8177, 25'd3217, 25'd13404, 25'd2681, 25'd17023}, '{25'd6032, 25'd10455, 25'd12466, 25'd1743, 25'd3619, -25'd4691, -25'd3619, 25'd7238, 25'd7640}, '{-25'd5362, -25'd10991, -25'd8311, -25'd2681, -25'd2547, -25'd938, 25'd12734, -25'd5496, 25'd11259}}, '{'{-25'd670, 25'd7506, 25'd4155, -25'd1877, -25'd6032, -25'd8981, -25'd1474, -25'd268, 25'd8445}, '{25'd0, 25'd4691, -25'd3083, -25'd2011, -25'd10187, 25'd5228, -25'd1072, -25'd5630, -25'd5630}, '{25'd6836, -25'd402, -25'd10321, -25'd5630, 25'd3887, -25'd7506, 25'd12466, -25'd6032, -25'd2279}, '{25'd268, 25'd11259, -25'd536, 25'd1206, -25'd7774, 25'd268, -25'd6970, 25'd3485, 25'd6836}, '{25'd9517, -25'd3217, 25'd2413, -25'd4423, -25'd938, 25'd6970, -25'd4691, -25'd8847, -25'd7908}, '{25'd10589, -25'd9517, 25'd7104, -25'd8177, -25'd7640, 25'd1474, -25'd3083, 25'd6032, 25'd7372}, '{-25'd4289, -25'd8981, 25'd9517, 25'd3753, -25'd3351, -25'd5094, 25'd1608, 25'd14610, 25'd10455}, '{25'd7238, -25'd134, 25'd804, 25'd1206, 25'd2547, -25'd402, -25'd1608, 25'd6434, -25'd6032}, '{25'd6300, 25'd5496, 25'd7104, 25'd5362, 25'd6434, 25'd11259, 25'd14879, 25'd13136, 25'd2547}}},
    '{'{'{25'd10454, -25'd3792, 25'd7892, -25'd1332, -25'd922, 25'd3075, 25'd5227, 25'd7379, -25'd10864}, '{-25'd4920, -25'd8917, -25'd9634, 25'd2460, 25'd9327, -25'd9942, -25'd3177, -25'd1947, -25'd4100}, '{25'd7789, 25'd1947, 25'd5125, 25'd9019, 25'd10762, 25'd11479, -25'd11069, -25'd2562, -25'd6149}, '{25'd1742, 25'd11274, -25'd1742, -25'd2460, 25'd8097, 25'd102, 25'd10762, -25'd3177, -25'd10454}, '{25'd7174, -25'd6867, 25'd10044, 25'd205, 25'd1845, -25'd1025, -25'd10557, -25'd5227, 25'd1435}, '{25'd9019, 25'd6252, -25'd4510, 25'd2767, -25'd102, 25'd10454, 25'd10762, -25'd7174, 25'd5842}, '{25'd3485, 25'd2562, 25'd5022, 25'd2562, 25'd10147, 25'd4612, -25'd10762, 25'd1640, 25'd1640}, '{-25'd7482, -25'd4920, 25'd10864, 25'd3792, 25'd12197, -25'd8302, 25'd4715, 25'd10864, -25'd5125}, '{25'd512, -25'd9942, -25'd3177, 25'd2562, 25'd6457, 25'd6252, -25'd9019, 25'd8917, -25'd4100}}, '{'{-25'd6559, 25'd6867, 25'd9737, 25'd6969, -25'd4305, -25'd5022, 25'd7072, -25'd5945, -25'd7379}, '{-25'd2255, -25'd4100, 25'd5330, 25'd10557, -25'd9224, -25'd10147, -25'd10044, 25'd7789, 25'd5842}, '{-25'd4100, -25'd922, 25'd0, 25'd7994, -25'd6867, -25'd5535, 25'd9942, 25'd4510, 25'd7277}, '{25'd8814, -25'd10557, -25'd2562, -25'd1742, 25'd0, 25'd6662, -25'd8507, -25'd10864, -25'd5740}, '{25'd6662, 25'd10044, 25'd10967, 25'd615, 25'd3177, -25'd11992, 25'd6252, -25'd9429, -25'd9019}, '{25'd5740, -25'd7687, 25'd7379, -25'd9532, -25'd10557, 25'd102, 25'd717, 25'd10454, 25'd10557}, '{25'd4407, 25'd9429, 25'd9942, 25'd2460, 25'd1435, 25'd4715, -25'd9839, 25'd5535, 25'd1435}, '{25'd1537, 25'd6354, 25'd1435, 25'd1640, -25'd11172, 25'd10454, -25'd10762, 25'd3280, 25'd5842}, '{-25'd11274, 25'd4920, 25'd3997, 25'd2357, 25'd8814, -25'd6559, 25'd9327, 25'd2562, 25'd6867}}, '{'{-25'd2562, -25'd10659, 25'd12299, 25'd9532, -25'd5330, -25'd5330, -25'd9839, 25'd11684, 25'd2460}, '{25'd6457, 25'd0, -25'd7379, -25'd7379, 25'd410, 25'd3690, -25'd1640, 25'd9532, -25'd2870}, '{25'd4510, -25'd6559, -25'd7482, -25'd410, 25'd3280, 25'd8609, -25'd2460, -25'd1435, 25'd9327}, '{25'd7994, 25'd10454, 25'd7277, 25'd5227, -25'd820, 25'd7892, -25'd205, -25'd6662, -25'd102}, '{25'd4305, 25'd3280, 25'd102, 25'd2460, -25'd5330, 25'd6457, 25'd8712, -25'd9737, 25'd2357}, '{-25'd7379, -25'd11172, 25'd1537, -25'd2050, 25'd10044, 25'd2460, 25'd4715, 25'd5535, 25'd13016}, '{-25'd4817, -25'd9839, 25'd10557, -25'd3792, 25'd3485, -25'd9019, -25'd3177, -25'd6252, -25'd717}, '{-25'd307, 25'd10864, 25'd2665, -25'd3485, -25'd9327, -25'd2562, 25'd1537, -25'd8609, 25'd512}, '{25'd3075, -25'd8814, 25'd10557, 25'd11684, 25'd3587, -25'd3792, -25'd9019, -25'd5330, 25'd7482}}},
    '{'{'{25'd11914, 25'd2383, -25'd2924, 25'd2058, 25'd4224, -25'd7474, -25'd8773, -25'd10073, 25'd9532}, '{25'd4657, 25'd4441, 25'd867, -25'd11048, 25'd4008, 25'd6932, -25'd10940, 25'd108, -25'd7149}, '{25'd650, -25'd7474, 25'd10723, 25'd10506, -25'd8448, 25'd2816, -25'd3791, 25'd9965, 25'd9315}, '{-25'd5091, 25'd2600, -25'd7040, -25'd7799, -25'd758, -25'd6932, -25'd10181, -25'd2058, -25'd5307}, '{25'd4008, -25'd1950, -25'd3683, -25'd10723, 25'd9532, -25'd10181, 25'd9423, 25'd4982, -25'd9098}, '{-25'd6282, -25'd2491, 25'd5524, -25'd1191, 25'd11806, 25'd8665, -25'd2383, 25'd1625, 25'd12131}, '{25'd9098, -25'd2924, 25'd108, -25'd2924, 25'd2708, 25'd4982, 25'd4549, 25'd12781, 25'd5416}, '{25'd8015, -25'd3141, 25'd3358, 25'd8124, -25'd8557, 25'd10615, -25'd1408, 25'd10073, 25'd8557}, '{25'd5632, -25'd5957, 25'd8448, -25'd3791, 25'd9315, 25'd3791, 25'd8773, -25'd4874, -25'd2275}}, '{'{25'd5416, -25'd13756, -25'd8990, -25'd1300, -25'd975, -25'd10181, -25'd9965, -25'd9532, 25'd7690}, '{-25'd7690, -25'd4224, -25'd3466, -25'd10181, -25'd6715, 25'd5632, -25'd650, 25'd8990, -25'd3358}, '{-25'd2058, -25'd8990, -25'd8665, -25'd12348, -25'd6066, 25'd2816, -25'd7365, 25'd1083, 25'd108}, '{-25'd6824, 25'd6282, -25'd2166, -25'd2708, 25'd542, 25'd4116, 25'd867, -25'd9748, -25'd4333}, '{-25'd3683, -25'd5416, -25'd1516, -25'd7690, -25'd4116, -25'd8340, 25'd7365, -25'd2708, -25'd9207}, '{25'd6174, 25'd9748, -25'd1191, 25'd3033, 25'd325, -25'd542, -25'd2924, -25'd6607, 25'd7365}, '{-25'd9965, 25'd5091, -25'd11806, -25'd325, -25'd3791, -25'd12348, -25'd12023, -25'd108, 25'd6066}, '{25'd6391, 25'd9532, -25'd1408, -25'd1083, -25'd8557, 25'd9640, -25'd8015, -25'd9423, 25'd9315}, '{-25'd11048, 25'd7582, 25'd2816, 25'd3249, -25'd2708, -25'd7365, -25'd12673, -25'd8557, 25'd3141}}, '{'{25'd5741, 25'd11914, -25'd1408, 25'd11481, 25'd2166, -25'd217, 25'd9857, -25'd8882, 25'd10615}, '{25'd3141, 25'd9965, 25'd758, -25'd975, 25'd5957, 25'd10831, 25'd8665, -25'd9640, 25'd12998}, '{-25'd9748, -25'd7582, 25'd2383, 25'd7582, 25'd1300, -25'd6066, 25'd1516, -25'd9207, 25'd1516}, '{25'd11914, -25'd3141, 25'd2275, 25'd5524, 25'd4874, 25'd10398, 25'd2383, 25'd9748, 25'd6824}, '{-25'd1516, -25'd1083, 25'd9423, -25'd11048, 25'd11373, -25'd1191, 25'd5957, 25'd3791, 25'd12889}, '{-25'd1733, -25'd5632, 25'd5741, 25'd2383, -25'd5741, 25'd217, 25'd433, 25'd1083, 25'd8773}, '{-25'd433, 25'd7907, 25'd758, -25'd975, -25'd975, 25'd0, 25'd5849, -25'd8015, -25'd7149}, '{-25'd6174, -25'd10073, -25'd542, 25'd8882, 25'd3249, 25'd5632, 25'd8665, 25'd12348, -25'd3249}, '{25'd2708, 25'd1408, -25'd9965, 25'd433, 25'd9207, -25'd6174, -25'd758, 25'd9965, 25'd8557}}},
    '{'{'{25'd3273, -25'd701, -25'd7481, -25'd2338, 25'd9702, -25'd12157, 25'd4676, 25'd4325, 25'd4208}, '{-25'd10520, 25'd11339, -25'd4091, -25'd6312, 25'd3156, -25'd4325, 25'd4208, -25'd4910, -25'd4910}, '{-25'd8650, 25'd1753, 25'd1637, 25'd5962, -25'd12040, 25'd468, 25'd5260, -25'd351, -25'd10754}, '{-25'd3273, -25'd6195, -25'd5728, -25'd10403, -25'd4208, 25'd6663, -25'd1286, -25'd1403, -25'd234}, '{-25'd8533, 25'd4793, 25'd117, -25'd11456, -25'd8299, 25'd8650, -25'd7481, -25'd8416, -25'd6546}, '{-25'd2338, 25'd468, 25'd7364, 25'd4325, 25'd3857, -25'd1637, 25'd3741, 25'd3156, -25'd8533}, '{25'd10520, -25'd9585, -25'd468, -25'd8066, 25'd8416, -25'd2805, -25'd8533, 25'd701, 25'd8183}, '{25'd6429, 25'd5962, 25'd3974, -25'd6546, 25'd5845, 25'd3741, -25'd1286, -25'd10637, -25'd10988}, '{-25'd10170, -25'd1286, -25'd2572, -25'd701, -25'd11572, -25'd8767, 25'd2805, -25'd9235, -25'd117}}, '{'{25'd3156, -25'd5260, -25'd8416, -25'd7832, 25'd3857, -25'd3507, -25'd6195, 25'd1637, 25'd4793}, '{25'd11105, -25'd2805, -25'd11923, -25'd3857, -25'd10637, 25'd351, -25'd1870, -25'd8066, -25'd9936}, '{25'd3507, -25'd1987, 25'd351, 25'd3039, 25'd5845, -25'd1753, 25'd5845, -25'd4559, 25'd1169}, '{-25'd3857, 25'd6195, 25'd3857, 25'd5845, -25'd4091, -25'd9702, -25'd9585, -25'd5260, -25'd4559}, '{-25'd12040, 25'd9001, -25'd10287, -25'd7949, -25'd818, 25'd8183, 25'd7014, 25'd9118, -25'd4793}, '{-25'd7832, 25'd10053, -25'd8533, 25'd8650, -25'd5728, -25'd6195, -25'd12858, -25'd7949, 25'd3273}, '{-25'd8533, 25'd8767, 25'd4208, 25'd3974, 25'd6897, -25'd935, 25'd10053, 25'd10053, -25'd8066}, '{25'd1403, -25'd7130, 25'd1637, -25'd6078, -25'd13326, -25'd9702, 25'd1286, -25'd11105, -25'd7364}, '{25'd9001, -25'd5962, -25'd12624, 25'd6780, -25'd468, 25'd3390, 25'd2689, -25'd1403, 25'd7949}}, '{'{-25'd2572, 25'd9351, 25'd14495, -25'd6312, 25'd13092, 25'd9936, 25'd6429, 25'd584, 25'd5377}, '{-25'd5845, 25'd1286, 25'd10403, 25'd8767, 25'd6429, 25'd13209, -25'd1520, -25'd7598, 25'd1403}, '{-25'd1870, -25'd6780, -25'd2221, 25'd8416, 25'd7715, 25'd4559, -25'd4208, 25'd4559, -25'd1520}, '{25'd2689, -25'd7598, 25'd13793, 25'd7247, 25'd3039, 25'd12391, -25'd4559, 25'd11806, -25'd818}, '{-25'd2455, 25'd7832, -25'd3974, -25'd3974, 25'd12040, 25'd701, 25'd11339, 25'd14845, 25'd5494}, '{25'd2572, 25'd8884, -25'd6429, -25'd5143, 25'd2455, 25'd9001, -25'd2572, -25'd7130, -25'd6312}, '{25'd11105, -25'd7715, -25'd4793, 25'd818, 25'd2805, 25'd11105, -25'd7949, 25'd9819, 25'd3039}, '{-25'd6897, 25'd1052, 25'd9235, 25'd584, 25'd2455, 25'd1169, 25'd11222, -25'd3273, -25'd3390}, '{25'd11339, 25'd12975, 25'd13209, -25'd3741, -25'd2572, -25'd2922, 25'd6078, -25'd6546, 25'd8884}}},
    '{'{'{25'd3009, 25'd7925, 25'd8627, 25'd8025, -25'd2608, 25'd3812, -25'd1003, 25'd7624, -25'd8025}, '{-25'd401, 25'd6320, -25'd1404, 25'd10132, -25'd502, 25'd7022, -25'd11335, -25'd7122, 25'd5016}, '{25'd3310, -25'd9329, 25'd3110, 25'd3310, 25'd10834, -25'd2809, 25'd1505, 25'd5617, 25'd5116}, '{-25'd7824, 25'd9329, 25'd702, 25'd7624, 25'd5718, 25'd903, 25'd10633, -25'd3812, 25'd6019}, '{-25'd702, -25'd903, 25'd4012, -25'd1103, -25'd6119, -25'd10432, 25'd8727, -25'd2809, 25'd4113}, '{-25'd12338, -25'd12138, -25'd8125, -25'd2407, 25'd8727, -25'd10232, 25'd5116, 25'd6821, 25'd3411}, '{25'd3812, 25'd6520, -25'd3310, 25'd6520, -25'd3812, -25'd6420, 25'd8226, -25'd1103, -25'd9931}, '{-25'd100, 25'd8326, 25'd10132, 25'd6119, -25'd9429, 25'd3812, -25'd6420, -25'd10031, -25'd10132}, '{-25'd4213, 25'd10834, -25'd2608, 25'd10934, -25'd5818, -25'd3511, -25'd11034, 25'd4715, -25'd11235}}, '{'{-25'd9028, 25'd7824, 25'd4414, -25'd11034, 25'd5317, 25'd4915, 25'd11436, -25'd7925, 25'd1705}, '{25'd4915, 25'd11536, -25'd4113, 25'd6621, -25'd9730, 25'd7724, 25'd201, -25'd7824, 25'd6019}, '{25'd1705, 25'd7122, -25'd7022, 25'd2708, 25'd8727, 25'd3812, 25'd2107, 25'd2809, 25'd7323}, '{-25'd9429, 25'd12740, 25'd2207, 25'd9730, 25'd6721, -25'd201, -25'd7323, -25'd10432, -25'd8827}, '{25'd6219, -25'd3712, -25'd4614, -25'd9831, 25'd5818, -25'd9630, 25'd7724, 25'd9730, 25'd10934}, '{-25'd2107, -25'd4414, -25'd3110, -25'd4012, 25'd10031, -25'd9229, 25'd2107, 25'd5216, -25'd9429}, '{-25'd1103, 25'd3210, -25'd8827, 25'd401, -25'd10633, -25'd3310, 25'd1705, -25'd4414, 25'd7624}, '{-25'd10834, -25'd8025, -25'd5216, 25'd2307, 25'd11034, 25'd11837, -25'd2107, -25'd5818, 25'd10132}, '{-25'd9931, -25'd7624, 25'd6922, 25'd10232, -25'd8326, 25'd3009, -25'd6420, -25'd9630, 25'd6019}}, '{'{-25'd6922, -25'd802, 25'd6420, 25'd11235, 25'd7624, 25'd4715, 25'd5918, 25'd4113, -25'd4815}, '{25'd10633, -25'd9028, -25'd6420, -25'd7925, 25'd502, -25'd4213, -25'd6420, 25'd903, 25'd2608}, '{25'd6721, 25'd3712, -25'd6119, -25'd5016, -25'd6621, 25'd7624, 25'd5517, -25'd2909, -25'd6520}, '{25'd11536, 25'd2307, 25'd6219, -25'd2809, -25'd6420, -25'd4614, 25'd7824, 25'd7423, 25'd9429}, '{-25'd2207, -25'd401, 25'd6922, 25'd7925, -25'd3009, 25'd3310, -25'd1204, -25'd4715, -25'd7624}, '{25'd3310, -25'd8727, 25'd10332, 25'd5317, 25'd3310, -25'd10031, 25'd7624, 25'd903, -25'd5016}, '{-25'd5016, 25'd12238, 25'd11135, 25'd6219, -25'd9931, -25'd2909, 25'd7523, -25'd3912, -25'd201}, '{-25'd401, -25'd10432, 25'd5016, -25'd3712, -25'd2107, -25'd8125, 25'd2207, -25'd3110, 25'd100}, '{25'd2107, -25'd6520, -25'd9630, -25'd502, -25'd8326, 25'd7624, 25'd11135, -25'd11636, 25'd7222}}},
    '{'{'{25'd5344, 25'd7391, -25'd9552, 25'd9893, -25'd8528, 25'd10803, 25'd12053, 25'd4435, 25'd11599}, '{-25'd455, 25'd12394, -25'd5003, 25'd1365, -25'd4662, 25'd12167, -25'd796, 25'd11599, -25'd1706}, '{25'd6823, 25'd11826, -25'd9552, -25'd3184, 25'd569, 25'd4776, -25'd9097, 25'd2502, -25'd1819}, '{25'd1251, 25'd1478, 25'd2274, 25'd12394, 25'd2274, -25'd569, 25'd12849, 25'd5117, -25'd3411}, '{25'd569, 25'd5003, -25'd7277, 25'd3298, 25'd2388, -25'd4094, -25'd7505, 25'd11030, -25'd5686}, '{-25'd6027, 25'd11485, 25'd910, 25'd5458, 25'd7050, 25'd7050, -25'd6254, -25'd7619, 25'd4094}, '{-25'd6254, 25'd4435, -25'd682, 25'd11371, 25'd2502, 25'd6254, -25'd1478, 25'd569, 25'd1819}, '{-25'd2274, 25'd13986, -25'd8301, -25'd8642, -25'd682, -25'd4435, -25'd7391, 25'd11257, -25'd8528}, '{25'd3980, -25'd569, 25'd7391, 25'd3411, 25'd3525, 25'd6027, 25'd2956, -25'd7732, -25'd6709}}, '{'{-25'd8756, -25'd10689, -25'd8301, -25'd10461, 25'd569, 25'd4321, -25'd7960, -25'd2047, -25'd6823}, '{-25'd8187, -25'd3298, 25'd1251, -25'd4321, 25'd4321, -25'd8983, -25'd13304, 25'd1819, -25'd3411}, '{-25'd10120, -25'd6482, 25'd3980, -25'd11144, 25'd114, 25'd8756, -25'd5003, 25'd569, 25'd5799}, '{25'd3639, 25'd6823, -25'd7960, 25'd8073, 25'd6368, -25'd13532, 25'd4321, -25'd12281, -25'd6368}, '{-25'd4435, 25'd1137, 25'd7050, -25'd7505, -25'd10348, -25'd341, -25'd10916, -25'd3298, -25'd5344}, '{-25'd10348, -25'd5344, -25'd5913, -25'd6595, -25'd910, 25'd455, -25'd14328, -25'd5799, -25'd4207}, '{-25'd13190, -25'd4776, 25'd7391, 25'd1478, -25'd4094, -25'd5913, -25'd7277, -25'd11485, 25'd1933}, '{-25'd6368, -25'd7619, -25'd1365, 25'd7050, -25'd1933, 25'd3980, 25'd2615, 25'd1023, 25'd5572}, '{-25'd6482, 25'd6368, -25'd682, -25'd1137, 25'd3752, -25'd2502, -25'd5003, -25'd10007, -25'd8415}}, '{'{-25'd1706, 25'd8073, -25'd5231, 25'd11485, 25'd7619, -25'd7505, -25'd3752, 25'd6140, -25'd10120}, '{25'd455, 25'd7164, -25'd5458, 25'd0, 25'd12167, 25'd8756, -25'd2161, 25'd1251, -25'd4776}, '{25'd11940, -25'd9211, 25'd5003, -25'd2274, 25'd12167, 25'd11599, 25'd9779, 25'd12167, -25'd1365}, '{25'd5458, 25'd9779, 25'd7050, -25'd1933, 25'd1933, -25'd1251, 25'd12167, 25'd9211, -25'd1706}, '{25'd6254, 25'd12167, 25'd5686, -25'd7619, 25'd1478, -25'd3298, 25'd227, -25'd10234, -25'd569}, '{25'd6709, -25'd4207, 25'd10916, -25'd5799, -25'd8073, -25'd5799, 25'd4776, -25'd2502, -25'd7050}, '{25'd10575, -25'd796, 25'd14441, 25'd5003, 25'd5117, 25'd11940, -25'd227, 25'd12736, 25'd6254}, '{25'd2274, 25'd796, 25'd6595, -25'd2047, 25'd1478, -25'd1365, -25'd3639, -25'd2274, 25'd1365}, '{25'd11371, 25'd682, 25'd1251, 25'd11144, -25'd3070, 25'd2502, 25'd11371, -25'd1365, 25'd4207}}},
    '{'{'{25'd5108, 25'd165, -25'd12357, 25'd2801, -25'd14829, -25'd2307, 25'd2142, 25'd1648, -25'd12687}, '{-25'd15982, -25'd13511, 25'd2636, -25'd6920, -25'd12687, -25'd11534, 25'd1648, 25'd2801, -25'd8897}, '{-25'd7414, -25'd16147, -25'd4449, -25'd15817, 25'd3295, -25'd824, -25'd12687, -25'd10710, -25'd13181}, '{-25'd1977, -25'd16971, -25'd7909, -25'd20596, 25'd1318, -25'd16147, 25'd4943, 25'd1153, -25'd5108}, '{-25'd13675, -25'd17300, -25'd16971, -25'd21090, -25'd8238, -25'd1812, -25'd1648, -25'd6261, -25'd4943}, '{25'd0, -25'd16147, -25'd8073, -25'd2966, -25'd5932, 25'd2307, -25'd13181, -25'd9062, -25'd9062}, '{-25'd13840, 25'd2142, -25'd16312, -25'd11863, -25'd3954, 25'd1318, 25'd8403, 25'd10051, 25'd4119}, '{-25'd2636, -25'd17136, -25'd5108, -25'd18124, -25'd17136, 25'd5108, 25'd8568, 25'd6920, -25'd1648}, '{-25'd3625, -25'd17136, -25'd6591, -25'd6426, -25'd6426, -25'd11534, -25'd1318, -25'd494, -25'd3460}}, '{'{25'd8238, 25'd2966, 25'd1318, 25'd2142, -25'd10545, 25'd0, 25'd9721, -25'd3131, 25'd6426}, '{25'd10874, 25'd6426, 25'd10545, 25'd2471, 25'd10215, 25'd10874, -25'd1977, -25'd8238, -25'd494}, '{25'd4119, 25'd3295, 25'd5767, -25'd4449, -25'd5272, -25'd659, 25'd1153, -25'd3460, 25'd9227}, '{25'd1977, -25'd7250, 25'd824, 25'd4613, -25'd3790, -25'd4449, 25'd1977, 25'd330, 25'd3295}, '{-25'd9227, -25'd4943, -25'd5932, -25'd2307, 25'd6426, 25'd11039, -25'd330, 25'd10215, 25'd6261}, '{25'd12522, 25'd1483, 25'd13016, 25'd7744, 25'd2142, 25'd11204, -25'd9392, -25'd989, -25'd330}, '{25'd10215, 25'd6426, 25'd1812, -25'd7744, 25'd3790, -25'd7744, -25'd3790, -25'd1153, 25'd2307}, '{-25'd8073, -25'd7579, 25'd5932, 25'd3460, -25'd2801, 25'd8568, 25'd4449, -25'd6920, 25'd2966}, '{25'd11204, 25'd659, 25'd5767, 25'd5272, 25'd6920, 25'd5437, 25'd6261, 25'd2636, -25'd1153}}, '{'{-25'd4119, -25'd7909, 25'd9392, 25'd7909, 25'd5602, 25'd1812, -25'd4449, 25'd8897, -25'd3790}, '{25'd659, 25'd1977, 25'd3625, 25'd2636, 25'd10874, -25'd4778, 25'd3954, -25'd5108, 25'd11698}, '{-25'd1483, 25'd3295, -25'd3790, 25'd1977, -25'd3954, 25'd7414, 25'd9392, 25'd7909, -25'd8073}, '{-25'd6755, -25'd4449, 25'd9556, 25'd11204, 25'd8403, -25'd9556, 25'd7579, 25'd10545, -25'd2966}, '{25'd8238, 25'd5272, -25'd9062, 25'd5767, -25'd8403, -25'd3131, 25'd494, 25'd4613, 25'd6261}, '{25'd9886, 25'd8238, -25'd5272, 25'd9556, 25'd11534, -25'd10380, -25'd6591, -25'd2471, -25'd9062}, '{25'd4284, 25'd2966, 25'd494, -25'd3460, -25'd4943, -25'd11039, 25'd9392, 25'd3131, -25'd6426}, '{-25'd7579, 25'd11039, 25'd5272, 25'd9886, 25'd7909, -25'd1483, -25'd4943, 25'd8897, -25'd9886}, '{-25'd3131, 25'd330, 25'd5272, -25'd659, 25'd3131, 25'd4943, -25'd7250, 25'd5932, 25'd4943}}},
    '{'{'{-25'd199, -25'd10134, 25'd7153, 25'd8147, -25'd8743, -25'd4769, 25'd5663, 25'd8644, 25'd2981}, '{-25'd298, -25'd6458, 25'd497, 25'd11128, 25'd3875, -25'd10333, 25'd5166, 25'd1987, 25'd5564}, '{25'd7849, -25'd1490, -25'd10830, -25'd5266, 25'd7551, 25'd2484, -25'd4272, 25'd4074, -25'd9836}, '{25'd2583, 25'd10233, 25'd3080, 25'd7452, 25'd3080, -25'd6557, 25'd199, 25'd10432, -25'd3875}, '{-25'd2484, 25'd8445, 25'd596, 25'd5365, -25'd7153, -25'd1292, 25'd2981, -25'd695, 25'd12618}, '{25'd7849, 25'd1391, 25'd1292, 25'd2285, 25'd2881, 25'd3676, -25'd2484, -25'd5365, 25'd12519}, '{-25'd5763, 25'd1490, 25'd11823, -25'd5663, -25'd2981, 25'd10532, -25'd6557, 25'd4670, -25'd7153}, '{25'd7750, 25'd9041, 25'd7352, -25'd894, -25'd2981, -25'd10333, 25'd11227, 25'd12121, -25'd8246}, '{-25'd4372, -25'd3477, 25'd1490, 25'd11426, 25'd2086, -25'd3378, -25'd5564, -25'd7153, -25'd1888}}, '{'{25'd3875, -25'd4670, 25'd11426, 25'd8445, -25'd2881, 25'd6955, -25'd8346, -25'd9439, -25'd3577}, '{25'd11624, 25'd2583, 25'd3775, 25'd596, 25'd7253, -25'd7551, -25'd1590, 25'd1292, 25'd2086}, '{25'd10830, 25'd10730, 25'd7551, 25'd2683, 25'd695, -25'd4769, 25'd4769, -25'd7352, -25'd7352}, '{25'd1093, -25'd2583, 25'd3775, -25'd596, 25'd9737, -25'd10432, 25'd9439, -25'd2086, -25'd10333}, '{-25'd2881, -25'd8743, -25'd9240, -25'd2186, -25'd5266, -25'd2186, -25'd5266, 25'd5266, -25'd8445}, '{-25'd6855, 25'd6359, 25'd5067, 25'd2086, 25'd9538, 25'd8445, -25'd8147, 25'd8743, 25'd9339}, '{25'd7750, 25'd1292, 25'd10830, 25'd7948, -25'd3378, -25'd7452, 25'd2285, -25'd2086, -25'd10532}, '{25'd12618, 25'd9439, -25'd8843, 25'd8644, 25'd1192, 25'd298, -25'd7253, -25'd397, -25'd10532}, '{25'd9439, 25'd11724, 25'd11326, -25'd8346, 25'd11823, -25'd8346, -25'd298, 25'd9041, -25'd3477}}, '{'{25'd8246, -25'd6458, -25'd10333, 25'd596, 25'd8644, -25'd298, -25'd695, -25'd3875, -25'd4670}, '{-25'd10532, 25'd3279, -25'd5763, 25'd5564, 25'd1590, -25'd9637, 25'd2981, -25'd4074, 25'd2285}, '{-25'd2086, 25'd1391, 25'd5564, -25'd4173, 25'd4769, 25'd11624, 25'd5564, -25'd11128, -25'd10035}, '{25'd3279, 25'd5961, 25'd9240, -25'd7253, 25'd2683, -25'd695, 25'd2981, 25'd10333, -25'd2583}, '{-25'd5067, -25'd1391, -25'd6756, 25'd5663, -25'd5166, -25'd7849, -25'd1888, 25'd894, 25'd4570}, '{25'd4372, -25'd9339, -25'd10035, -25'd7551, -25'd795, -25'd4471, -25'd10333, 25'd9538, 25'd1192}, '{25'd6955, 25'd10830, -25'd9538, 25'd4868, -25'd5067, 25'd1788, -25'd1987, -25'd9836, -25'd6955}, '{25'd3676, -25'd7054, -25'd7750, 25'd3378, 25'd11128, 25'd3378, 25'd2086, 25'd1192, 25'd5862}, '{-25'd7452, -25'd1987, 25'd8048, 25'd8942, 25'd9339, -25'd11227, 25'd9538, 25'd11326, -25'd11326}}},
    '{'{'{25'd11464, -25'd4425, -25'd2916, -25'd6034, 25'd8045, 25'd402, -25'd6235, 25'd4927, 25'd12771}, '{25'd603, 25'd3117, 25'd8246, 25'd5832, 25'd12168, 25'd10961, -25'd6436, 25'd8548, 25'd9252}, '{25'd4324, 25'd9654, 25'd8548, 25'd8950, 25'd0, -25'd8749, 25'd7341, -25'd8950, 25'd11665}, '{-25'd2615, 25'd2413, 25'd3520, -25'd2816, 25'd101, 25'd2916, 25'd10358, -25'd7844, -25'd8145}, '{25'd704, 25'd7039, 25'd603, -25'd10056, 25'd5430, -25'd7341, -25'd3620, -25'd10056, -25'd6134}, '{25'd2413, 25'd7441, -25'd10961, 25'd10559, 25'd5631, 25'd12570, -25'd10861, -25'd1810, 25'd2212}, '{-25'd8447, 25'd5330, -25'd1810, -25'd8950, 25'd12369, -25'd3419, 25'd6738, -25'd5229, 25'd3721}, '{25'd10861, -25'd9553, -25'd7039, 25'd5229, 25'd8347, 25'd12268, -25'd8246, -25'd2112, 25'd1307}, '{25'd9252, -25'd4425, -25'd6134, 25'd4626, 25'd6838, -25'd3821, 25'd9754, 25'd8648, 25'd8045}}, '{'{25'd8749, 25'd2212, -25'd6637, 25'd6738, 25'd4626, -25'd4525, 25'd8045, -25'd10257, 25'd11263}, '{-25'd9654, -25'd11766, 25'd5933, 25'd5832, -25'd11464, -25'd11464, 25'd9252, 25'd10458, 25'd6436}, '{25'd10056, 25'd201, -25'd9654, -25'd603, -25'd11162, -25'd4525, 25'd9553, 25'd8849, 25'd11766}, '{-25'd10157, -25'd6838, -25'd7643, 25'd5229, -25'd10861, -25'd5229, -25'd7039, -25'd11062, 25'd10257}, '{-25'd704, 25'd3620, 25'd503, -25'd8950, -25'd2715, 25'd11464, -25'd7643, 25'd603, 25'd11564}, '{25'd2615, -25'd1408, -25'd1810, 25'd7039, 25'd3821, -25'd9050, -25'd804, 25'd4324, -25'd7844}, '{25'd7643, -25'd6939, -25'd5330, -25'd7441, 25'd5933, 25'd6134, 25'd10458, 25'd7542, -25'd1508}, '{-25'd11162, -25'd101, 25'd6134, -25'd2816, -25'd1207, -25'd4224, -25'd3922, 25'd5832, 25'd6034}, '{25'd1710, 25'd2715, 25'd704, 25'd9050, -25'd9151, 25'd7944, -25'd9955, 25'd7441, 25'd2112}}, '{'{-25'd8849, 25'd11363, 25'd6335, 25'd11062, -25'd4827, -25'd804, 25'd9754, -25'd8648, -25'd10257}, '{25'd10659, 25'd11363, -25'd5531, 25'd1911, 25'd6939, 25'd7441, -25'd5531, 25'd7341, -25'd5933}, '{25'd6536, -25'd5330, -25'd7643, 25'd11665, -25'd4726, -25'd10257, 25'd10961, 25'd2715, -25'd3821}, '{25'd2916, -25'd603, -25'd1408, -25'd4123, -25'd3721, 25'd503, -25'd10157, -25'd1508, -25'd1609}, '{25'd1911, 25'd7844, -25'd10458, 25'd11866, 25'd10760, 25'd6235, 25'd7542, -25'd10659, 25'd3218}, '{25'd6034, 25'd5430, 25'd2816, -25'd9453, 25'd9855, -25'd3318, 25'd1307, 25'd11967, 25'd603}, '{-25'd1508, 25'd4927, -25'd3117, -25'd6235, -25'd4827, -25'd7039, 25'd2916, 25'd9754, 25'd1106}, '{25'd11162, 25'd8950, -25'd1106, -25'd6034, -25'd4525, 25'd10559, -25'd9352, 25'd6034, 25'd12570}, '{-25'd4726, -25'd8548, 25'd7441, -25'd10257, -25'd8246, 25'd4022, 25'd1508, 25'd10257, -25'd804}}},
    '{'{'{25'd6787, 25'd392, -25'd4046, 25'd12400, 25'd9006, -25'd1044, -25'd2611, -25'd6004, -25'd2350}, '{25'd4568, 25'd5091, 25'd522, -25'd783, 25'd5874, 25'd3133, 25'd5352, 25'd9529, 25'd783}, '{-25'd6135, 25'd5874, -25'd8484, -25'd8484, 25'd4046, 25'd4438, -25'd12270, -25'd9529, 25'd10181}, '{-25'd5743, -25'd1697, 25'd10573, 25'd6657, -25'd1436, -25'd10051, -25'd1305, 25'd5352, -25'd2480}, '{-25'd9659, 25'd10964, 25'd4307, 25'd8354, -25'd6396, 25'd5091, 25'd7310, -25'd5874, 25'd8615}, '{-25'd6004, 25'd3002, -25'd1305, 25'd4046, -25'd131, -25'd8484, 25'd3394, 25'd11356, -25'd4438}, '{-25'd5482, 25'd8354, -25'd6526, 25'd14489, -25'd5482, -25'd6396, -25'd5482, -25'd783, -25'd1436}, '{25'd7571, 25'd1958, -25'd1566, 25'd6657, -25'd7571, -25'd9529, 25'd7310, -25'd914, -25'd1958}, '{25'd3002, 25'd4438, 25'd11748, 25'd3263, -25'd6135, 25'd11748, -25'd5221, 25'd5091, 25'd4307}}, '{'{25'd11356, 25'd9006, 25'd8745, 25'd10834, -25'd7962, 25'd4699, -25'd3524, 25'd9137, -25'd13053}, '{-25'd9920, -25'd4046, 25'd11095, 25'd5352, 25'd13053, -25'd11748, -25'd12922, -25'd8223, 25'd1436}, '{25'd7310, 25'd9790, 25'd1566, -25'd5091, 25'd2350, -25'd6396, -25'd5221, 25'd7440, 25'd1566}, '{25'd9137, -25'd1566, 25'd1958, -25'd5091, -25'd8354, 25'd3394, -25'd7962, 25'd1697, -25'd12792}, '{-25'd7440, -25'd5091, 25'd1305, 25'd7179, 25'd1044, -25'd7962, -25'd12270, -25'd10834, -25'd4960}, '{-25'd8223, -25'd8223, -25'd9790, 25'd9659, -25'd783, -25'd7179, -25'd8484, -25'd7571, -25'd4568}, '{25'd8484, 25'd3002, 25'd5091, -25'd653, 25'd10051, 25'd914, 25'd5221, 25'd2219, -25'd13575}, '{-25'd8745, -25'd653, 25'd4046, 25'd3655, -25'd1566, -25'd7962, 25'd6918, 25'd5352, 25'd3785}, '{25'd1697, -25'd6004, 25'd11486, -25'd261, -25'd6657, -25'd8354, -25'd8615, -25'd9790, 25'd6787}}, '{'{25'd392, 25'd11356, 25'd1436, 25'd9659, 25'd13183, -25'd5352, 25'd2350, -25'd3524, -25'd914}, '{-25'd6265, 25'd12009, 25'd12270, -25'd2219, 25'd15272, -25'd3133, 25'd8484, -25'd4177, 25'd9659}, '{-25'd1305, 25'd1566, -25'd6004, 25'd9920, 25'd6787, -25'd3394, -25'd2741, -25'd1044, 25'd5482}, '{25'd9529, 25'd10442, 25'd14489, -25'd4830, 25'd7962, -25'd8484, 25'd13444, 25'd3916, 25'd10834}, '{25'd9659, 25'd12661, -25'd5482, 25'd12270, 25'd4438, -25'd8354, 25'd653, -25'd4046, 25'd9920}, '{-25'd4177, 25'd4960, 25'd5613, -25'd2611, -25'd2741, 25'd8615, 25'd1958, 25'd12792, 25'd3655}, '{25'd8484, -25'd4960, 25'd9398, 25'd11878, 25'd16055, -25'd8223, -25'd3916, 25'd5874, 25'd1044}, '{25'd5743, -25'd4830, 25'd16577, -25'd3655, 25'd2088, -25'd7962, -25'd5482, 25'd2350, 25'd0}, '{-25'd3263, 25'd13053, -25'd6657, -25'd6004, 25'd1175, 25'd11095, 25'd10181, 25'd15272, 25'd653}}},
    '{'{'{-25'd13005, -25'd9139, -25'd6327, 25'd2578, 25'd4921, -25'd6444, -25'd1757, -25'd9373, -25'd117}, '{25'd9022, -25'd11833, 25'd3398, -25'd8201, -25'd2929, -25'd6913, 25'd12068, 25'd9490, -25'd11013}, '{25'd2578, -25'd5389, -25'd13239, -25'd1523, 25'd10662, 25'd7030, -25'd11130, 25'd8553, -25'd11130}, '{-25'd1172, -25'd8436, 25'd7264, -25'd2578, 25'd5507, -25'd10779, -25'd586, -25'd10896, 25'd117}, '{25'd5507, 25'd9959, -25'd4218, -25'd4335, -25'd1992, -25'd6327, -25'd2695, 25'd8436, 25'd3281}, '{-25'd12302, 25'd5624, -25'd7967, -25'd9842, 25'd10779, 25'd1875, 25'd9022, 25'd9139, 25'd7264}, '{-25'd3749, -25'd8201, 25'd10310, -25'd8319, -25'd8201, 25'd3281, 25'd9607, -25'd6678, -25'd11716}, '{-25'd6210, 25'd351, 25'd469, 25'd6913, 25'd8319, 25'd2812, -25'd13357, -25'd11365, -25'd9959}, '{-25'd11013, -25'd234, 25'd1406, -25'd13239, -25'd6795, -25'd11833, -25'd11833, -25'd14060, -25'd14997}}, '{'{25'd10076, -25'd4452, -25'd7616, -25'd8553, 25'd10779, -25'd6561, 25'd2578, -25'd9607, -25'd2695}, '{-25'd5975, -25'd7264, -25'd6210, -25'd2226, 25'd12068, -25'd9490, 25'd7381, -25'd10193, -25'd937}, '{25'd7498, -25'd937, 25'd9256, -25'd6678, 25'd8553, 25'd12185, -25'd7850, 25'd8319, -25'd703}, '{-25'd10193, 25'd9842, -25'd2695, 25'd4101, -25'd937, -25'd820, 25'd12654, -25'd4687, 25'd3398}, '{-25'd7264, -25'd2460, 25'd6444, -25'd3749, 25'd4569, 25'd4335, 25'd2812, -25'd5155, 25'd12419}, '{25'd8319, -25'd5624, 25'd12536, -25'd2460, 25'd3163, 25'd9373, 25'd10076, -25'd1054, -25'd3866}, '{25'd117, 25'd4687, 25'd10076, 25'd6913, -25'd5038, -25'd9022, 25'd9022, -25'd8201, 25'd7498}, '{25'd1406, -25'd6913, 25'd12302, 25'd6795, -25'd820, 25'd4921, 25'd13122, -25'd2343, 25'd5272}, '{-25'd937, 25'd12771, 25'd10896, 25'd9842, 25'd13122, -25'd4218, 25'd9022, 25'd4921, 25'd234}}, '{'{25'd1875, 25'd2812, 25'd7616, -25'd5975, 25'd9256, -25'd6795, -25'd5975, 25'd12302, -25'd4569}, '{25'd11951, 25'd7147, -25'd9022, 25'd2226, -25'd2929, -25'd6561, 25'd1992, 25'd10427, 25'd5038}, '{25'd11248, -25'd8553, 25'd5507, 25'd10545, -25'd2812, -25'd2460, 25'd234, 25'd8787, 25'd3632}, '{25'd3515, 25'd2460, -25'd586, -25'd6795, 25'd6444, -25'd9607, 25'd469, -25'd11130, 25'd3398}, '{25'd7147, 25'd11833, 25'd2460, -25'd6092, 25'd8670, -25'd6561, 25'd11248, -25'd3046, -25'd117}, '{25'd10662, -25'd3163, -25'd11130, -25'd1875, -25'd4687, -25'd7616, -25'd7030, 25'd6444, 25'd8787}, '{25'd2578, -25'd9256, -25'd2812, 25'd6678, 25'd1406, 25'd7733, -25'd2695, 25'd9022, 25'd5272}, '{-25'd703, -25'd1289, -25'd6444, -25'd9373, -25'd9373, -25'd6327, 25'd7733, -25'd10662, 25'd2812}, '{-25'd6561, -25'd4687, -25'd1757, 25'd11130, 25'd7498, -25'd7381, -25'd4569, 25'd7030, 25'd8436}}},
    '{'{'{25'd4090, 25'd8540, 25'd7939, 25'd1203, 25'd12148, -25'd3729, 25'd6736, 25'd15276, 25'd9863}, '{25'd10825, 25'd3488, -25'd7578, 25'd13592, 25'd5172, 25'd8660, 25'd12389, 25'd8179, -25'd1804}, '{-25'd6615, -25'd9863, -25'd3729, 25'd6856, -25'd9021, 25'd2526, 25'd3608, 25'd9983, 25'd9262}, '{25'd7337, -25'd3729, -25'd5292, 25'd7578, 25'd10946, 25'd12629, 25'd6255, -25'd481, 25'd1083}, '{25'd1564, 25'd1323, -25'd8179, -25'd2285, 25'd9743, 25'd8901, -25'd10224, -25'd5052, -25'd5413}, '{-25'd10825, 25'd6134, -25'd4811, -25'd8901, -25'd5172, -25'd6255, -25'd9262, 25'd4450, -25'd8059}, '{-25'd7939, 25'd5653, -25'd10224, 25'd1203, 25'd9502, 25'd5052, 25'd2887, -25'd9863, 25'd6736}, '{-25'd6495, -25'd4811, -25'd10104, -25'd3849, -25'd1684, -25'd1443, -25'd3127, 25'd1323, -25'd6134}, '{-25'd9262, 25'd11186, 25'd4811, 25'd12990, -25'd10224, 25'd1323, -25'd8299, -25'd7097, -25'd120}}, '{'{-25'd7939, -25'd4090, -25'd120, -25'd10825, 25'd2045, -25'd1924, 25'd2045, 25'd4932, -25'd6014}, '{-25'd6495, -25'd5773, -25'd3368, 25'd8420, 25'd1924, 25'd8901, 25'd4090, 25'd7457, 25'd11908}, '{25'd1924, -25'd1924, -25'd10585, -25'd3368, 25'd7097, -25'd8179, 25'd3849, -25'd10344, -25'd4330}, '{25'd722, 25'd10344, -25'd3729, 25'd842, 25'd8059, -25'd9021, -25'd9863, -25'd722, -25'd8299}, '{25'd4571, 25'd11547, 25'd0, -25'd6014, -25'd7337, -25'd12750, 25'd9983, -25'd3007, -25'd12389}, '{-25'd9863, -25'd8059, 25'd6615, -25'd11908, -25'd5894, -25'd4450, -25'd1443, 25'd2406, -25'd241}, '{25'd5172, -25'd361, 25'd10464, -25'd1323, 25'd3248, -25'd962, -25'd7217, 25'd9262, -25'd9141}, '{-25'd2406, -25'd5172, -25'd1203, 25'd6014, -25'd1804, 25'd10344, -25'd4450, -25'd9382, 25'd4090}, '{-25'd9983, -25'd5653, -25'd8540, 25'd4932, -25'd4932, 25'd6615, 25'd2526, -25'd10825, -25'd4691}}, '{'{25'd11547, -25'd120, 25'd3127, -25'd3729, 25'd2766, -25'd3248, -25'd5172, -25'd9141, 25'd2045}, '{25'd3608, -25'd2526, 25'd5533, -25'd7578, 25'd1804, -25'd120, -25'd6495, 25'd5533, 25'd11306}, '{-25'd1083, 25'd120, -25'd8540, 25'd4571, 25'd962, -25'd5172, 25'd9502, 25'd7939, 25'd4571}, '{25'd6495, 25'd9262, 25'd9262, -25'd4210, -25'd2526, 25'd5172, 25'd8299, 25'd9502, 25'd1804}, '{-25'd7818, 25'd10946, 25'd12028, 25'd481, -25'd9622, 25'd3368, 25'd3849, -25'd8901, -25'd1804}, '{25'd7217, 25'd4691, 25'd4450, -25'd9141, 25'd12389, -25'd7578, -25'd3488, 25'd12629, 25'd2045}, '{25'd2646, -25'd9743, 25'd9502, -25'd6736, 25'd5172, -25'd1924, 25'd5172, 25'd10344, 25'd5653}, '{-25'd7217, 25'd601, -25'd1443, -25'd3248, 25'd10585, -25'd7337, 25'd5172, -25'd3248, -25'd2646}, '{25'd6736, 25'd4571, 25'd4811, -25'd241, 25'd1684, -25'd6255, -25'd5653, 25'd9983, -25'd1323}}},
    '{'{'{-25'd11111, -25'd10678, 25'd1010, -25'd9091, -25'd2597, -25'd11977, -25'd14430, -25'd18326, -25'd17460}, '{-25'd11255, 25'd4185, -25'd10245, -25'd866, 25'd8514, 25'd10390, -25'd17605, -25'd10245, 25'd577}, '{-25'd4329, -25'd3463, -25'd4618, 25'd144, 25'd4185, 25'd10967, 25'd722, -25'd6494, -25'd3608}, '{25'd6349, -25'd4040, 25'd5628, 25'd7215, 25'd8802, 25'd2309, 25'd3896, -25'd3463, 25'd8802}, '{25'd10823, 25'd9812, -25'd10534, -25'd6205, -25'd8081, 25'd2453, -25'd7359, -25'd11688, 25'd4040}, '{25'd11111, 25'd3752, -25'd5628, -25'd577, 25'd6349, -25'd1154, -25'd12699, 25'd9524, 25'd8658}, '{25'd1443, 25'd8225, -25'd1732, 25'd8225, 25'd9091, 25'd2020, 25'd11400, -25'd2165, 25'd12410}, '{-25'd7071, 25'd4762, -25'd6205, 25'd5483, -25'd7359, 25'd1443, -25'd12121, 25'd7071, 25'd3319}, '{-25'd866, -25'd7504, -25'd9235, 25'd8658, 25'd5628, -25'd5339, -25'd7215, -25'd12987, -25'd9524}}, '{'{25'd2453, -25'd3175, -25'd15296, 25'd9091, 25'd6494, 25'd16017, -25'd8225, -25'd4040, 25'd7215}, '{-25'd9668, 25'd2742, -25'd722, 25'd7071, -25'd4185, -25'd3030, 25'd9380, -25'd3175, 25'd4906}, '{-25'd1732, -25'd2742, -25'd3319, -25'd6926, -25'd2742, 25'd722, -25'd3608, -25'd3752, 25'd12843}, '{-25'd5483, 25'd7215, 25'd577, 25'd3752, -25'd8947, -25'd2742, 25'd4906, 25'd8081, 25'd3030}, '{-25'd1154, 25'd5339, -25'd1154, -25'd13997, 25'd3030, -25'd6638, -25'd8514, 25'd7359, 25'd4040}, '{25'd5916, -25'd10967, 25'd6494, -25'd10390, -25'd7504, 25'd6494, -25'd2742, -25'd10534, -25'd4762}, '{-25'd5195, -25'd15007, -25'd12266, -25'd10245, -25'd9091, 25'd11400, 25'd6349, 25'd6494, -25'd9668}, '{-25'd9091, -25'd6349, -25'd12699, -25'd433, 25'd4329, -25'd7937, 25'd3175, -25'd2020, 25'd4473}, '{-25'd4185, -25'd4906, -25'd4762, -25'd16306, 25'd5916, -25'd7359, -25'd2165, -25'd7504, 25'd2309}}, '{'{25'd8369, -25'd433, 25'd2597, -25'd13420, -25'd10390, -25'd6782, -25'd12843, -25'd18038, -25'd14430}, '{-25'd2020, -25'd144, -25'd6638, -25'd289, 25'd9957, -25'd15152, 25'd144, -25'd8081, -25'd8081}, '{25'd9812, 25'd7359, 25'd6205, 25'd2742, 25'd2886, -25'd3175, -25'd4185, -25'd12266, 25'd3319}, '{25'd12843, -25'd3030, -25'd2742, 25'd8514, 25'd2020, 25'd2453, 25'd3175, 25'd10101, 25'd10967}, '{-25'd1154, 25'd1299, -25'd5051, 25'd1587, -25'd4473, 25'd12843, 25'd5628, -25'd866, -25'd6782}, '{25'd14286, 25'd7071, 25'd7648, 25'd12843, -25'd4762, 25'd8947, -25'd9957, 25'd11255, 25'd3896}, '{-25'd1299, -25'd2165, -25'd4185, 25'd5339, -25'd2453, -25'd4040, -25'd11688, -25'd8947, -25'd3896}, '{-25'd7504, -25'd3175, 25'd4185, 25'd5483, -25'd4040, -25'd6926, -25'd12699, -25'd9524, -25'd9091}, '{25'd12266, 25'd6494, -25'd7792, 25'd7359, -25'd8081, -25'd3175, 25'd4473, -25'd9091, -25'd7215}}},
    '{'{'{-25'd5802, 25'd7403, 25'd1401, -25'd800, -25'd1701, 25'd5502, 25'd9704, -25'd3001, 25'd4802}, '{-25'd4902, 25'd3301, 25'd7703, 25'd10404, -25'd11004, 25'd900, -25'd6302, 25'd100, 25'd8503}, '{-25'd3001, -25'd8403, 25'd2801, -25'd7603, -25'd6402, -25'd2501, -25'd4502, -25'd1701, 25'd12705}, '{-25'd10004, 25'd1000, 25'd9504, -25'd7203, 25'd1901, 25'd6102, -25'd400, 25'd10904, -25'd10704}, '{-25'd9904, 25'd7203, 25'd7503, -25'd1200, -25'd100, 25'd11804, 25'd7903, 25'd11004, -25'd900}, '{25'd12705, 25'd3401, -25'd3901, -25'd6903, -25'd2801, 25'd10204, 25'd5402, 25'd11804, 25'd8003}, '{25'd5702, -25'd1801, -25'd5502, 25'd6402, 25'd11604, 25'd12305, 25'd12705, 25'd10704, -25'd1000}, '{25'd0, 25'd6102, -25'd8503, 25'd2401, -25'd11204, -25'd2001, 25'd6502, -25'd2301, -25'd3601}, '{-25'd5902, 25'd9203, -25'd4402, 25'd8903, -25'd1200, 25'd10104, -25'd8103, -25'd3501, 25'd11604}}, '{'{-25'd3901, -25'd10604, -25'd8803, 25'd1401, 25'd900, -25'd9303, 25'd6302, -25'd8103, -25'd200}, '{-25'd8303, -25'd9003, -25'd1501, -25'd7303, 25'd4602, 25'd11404, -25'd8203, 25'd11904, 25'd9804}, '{25'd2601, 25'd8603, -25'd6602, 25'd6502, 25'd4902, -25'd200, 25'd4102, -25'd9504, -25'd6502}, '{-25'd7303, 25'd11404, -25'd700, -25'd7603, 25'd11004, 25'd5502, 25'd3601, 25'd8203, 25'd1901}, '{25'd4702, 25'd5702, 25'd4802, 25'd7303, 25'd12005, -25'd1401, -25'd6302, 25'd4202, 25'd5702}, '{-25'd4102, -25'd1601, -25'd1701, 25'd1000, 25'd9604, -25'd8103, -25'd6202, -25'd8703, 25'd8703}, '{25'd1601, 25'd1000, -25'd8603, 25'd3501, 25'd6202, 25'd8603, 25'd4102, -25'd10204, -25'd6903}, '{25'd400, 25'd12205, 25'd4902, 25'd4402, 25'd800, -25'd7603, 25'd8803, 25'd5002, 25'd11204}, '{25'd800, -25'd4202, -25'd6002, -25'd300, 25'd6602, 25'd12105, 25'd1200, 25'd8303, 25'd9704}}, '{'{25'd11104, 25'd700, 25'd7703, 25'd7003, -25'd5902, -25'd7503, 25'd5802, 25'd2601, 25'd6703}, '{25'd700, 25'd2901, 25'd9604, -25'd5502, -25'd1000, 25'd8903, 25'd9003, 25'd2501, 25'd2501}, '{-25'd700, 25'd7003, -25'd600, 25'd3101, -25'd11804, -25'd10104, -25'd3001, -25'd4102, -25'd2701}, '{-25'd600, 25'd5802, -25'd500, -25'd8703, 25'd5002, -25'd6903, -25'd9804, -25'd1100, -25'd8303}, '{-25'd2501, 25'd9504, 25'd7003, 25'd4802, -25'd6502, -25'd9604, 25'd900, 25'd7903, 25'd6402}, '{25'd5302, 25'd8403, 25'd1501, -25'd9704, 25'd9504, -25'd4802, 25'd8703, -25'd1000, 25'd6703}, '{-25'd4602, 25'd5402, 25'd10404, 25'd6402, 25'd10304, -25'd10504, 25'd2101, 25'd9804, -25'd300}, '{25'd11104, 25'd7103, 25'd2001, -25'd500, -25'd9404, -25'd3601, -25'd6202, -25'd5302, 25'd700}, '{-25'd10104, -25'd3101, 25'd10904, -25'd4802, -25'd3601, 25'd10204, 25'd2601, -25'd8603, 25'd6502}}},
    '{'{'{-25'd6000, 25'd9530, -25'd5530, 25'd6942, 25'd4941, 25'd9765, 25'd4000, 25'd9295, -25'd2706}, '{25'd5412, -25'd1529, 25'd6706, 25'd4353, 25'd5412, 25'd4236, 25'd7177, 25'd1647, -25'd3412}, '{25'd3412, -25'd10354, 25'd11059, 25'd2706, -25'd12471, -25'd3294, -25'd5294, 25'd7177, -25'd4236}, '{25'd6942, -25'd2353, -25'd941, -25'd1177, -25'd7412, -25'd5765, 25'd3412, -25'd4000, -25'd1412}, '{-25'd10236, -25'd2000, 25'd1294, 25'd2353, -25'd11530, -25'd9648, -25'd7883, -25'd3530, 25'd2235}, '{25'd11295, -25'd11412, -25'd1765, -25'd5765, -25'd6824, -25'd2118, 25'd2235, 25'd6471, -25'd1529}, '{-25'd706, -25'd10236, -25'd6706, 25'd1529, -25'd8824, 25'd8118, -25'd5294, 25'd2353, 25'd7412}, '{25'd5530, -25'd1765, -25'd3412, 25'd8118, 25'd5883, 25'd9177, 25'd6353, -25'd2235, 25'd2353}, '{-25'd1765, -25'd1765, -25'd11648, -25'd7177, 25'd3530, 25'd3883, 25'd10589, 25'd941, 25'd1765}}, '{'{-25'd3412, -25'd9177, -25'd9648, -25'd9412, 25'd8000, 25'd353, -25'd3530, 25'd11177, 25'd8471}, '{-25'd6824, -25'd824, 25'd8589, -25'd7765, 25'd471, -25'd6236, 25'd4236, 25'd12001, 25'd824}, '{-25'd9412, 25'd8118, 25'd11177, 25'd1294, -25'd8942, 25'd11295, 25'd4588, 25'd11295, 25'd10354}, '{-25'd1529, -25'd11177, 25'd4353, 25'd2706, 25'd4824, 25'd588, -25'd2118, 25'd7295, -25'd9765}, '{25'd2235, 25'd1294, 25'd9177, -25'd10942, -25'd3412, 25'd2235, -25'd2000, -25'd4941, 25'd3059}, '{25'd3412, -25'd3530, 25'd8706, 25'd11765, 25'd8353, -25'd6000, 25'd5059, 25'd2941, 25'd5530}, '{-25'd7647, 25'd0, 25'd11530, -25'd5765, -25'd4706, -25'd4353, 25'd6353, 25'd9177, 25'd14942}, '{-25'd5647, 25'd2353, -25'd5883, -25'd2471, 25'd4471, -25'd6706, 25'd1294, 25'd2824, 25'd2353}, '{25'd8118, -25'd3177, -25'd1177, 25'd4118, -25'd8353, 25'd8589, -25'd8706, 25'd10118, 25'd2000}}, '{'{25'd2588, 25'd4824, 25'd11765, -25'd3294, -25'd10354, 25'd7530, 25'd706, -25'd4000, -25'd11177}, '{-25'd10706, 25'd10471, 25'd11530, 25'd1294, -25'd6824, -25'd5177, 25'd471, -25'd3059, 25'd3883}, '{25'd2000, 25'd8353, -25'd4000, 25'd10706, -25'd7295, 25'd7412, 25'd9883, 25'd2706, -25'd4706}, '{-25'd4941, 25'd10824, 25'd6706, -25'd4588, -25'd6353, 25'd3059, -25'd2471, 25'd5177, 25'd9765}, '{25'd4941, 25'd11059, -25'd1412, 25'd2000, -25'd3412, -25'd6942, -25'd1059, 25'd6471, -25'd5883}, '{25'd941, 25'd8706, -25'd9177, -25'd2588, 25'd588, -25'd2471, -25'd11295, -25'd10706, -25'd6824}, '{-25'd9530, 25'd8236, 25'd7765, 25'd6353, -25'd3177, 25'd5412, -25'd5765, -25'd7059, -25'd10001}, '{-25'd7177, -25'd5177, 25'd588, 25'd8236, -25'd7647, 25'd8471, -25'd8824, 25'd5412, 25'd1059}, '{25'd9530, 25'd4236, -25'd353, 25'd4118, -25'd10001, 25'd8942, -25'd8236, -25'd2471, -25'd5883}}},
    '{'{'{-25'd5247, -25'd9619, -25'd3716, 25'd8307, 25'd7542, 25'd8416, 25'd4809, 25'd1967, 25'd4700}, '{25'd9072, 25'd7979, 25'd10930, 25'd547, 25'd6558, -25'd10930, -25'd4919, 25'd4263, -25'd7651}, '{-25'd2077, -25'd765, -25'd10821, -25'd7761, -25'd10275, 25'd656, -25'd5793, 25'd9072, 25'd8416}, '{-25'd4263, 25'd5793, 25'd9291, 25'd9728, 25'd874, 25'd11368, 25'd3607, 25'd4809, 25'd3716}, '{25'd1749, 25'd6886, 25'd1093, 25'd1967, -25'd1967, 25'd10603, -25'd7870, -25'd2842, 25'd7761}, '{25'd4372, 25'd6121, 25'd4481, 25'd5575, -25'd2951, 25'd12351, -25'd328, -25'd4263, -25'd8854}, '{-25'd5247, 25'd8089, 25'd8526, 25'd7105, -25'd7870, 25'd8198, 25'd9072, -25'd874, 25'd4591}, '{25'd5793, 25'd7105, -25'd3498, -25'd4372, 25'd328, 25'd11149, 25'd1312, -25'd4263, 25'd12679}, '{-25'd7433, 25'd7214, 25'd765, 25'd4154, 25'd4154, -25'd656, 25'd1749, -25'd2951, 25'd5028}}, '{'{-25'd6230, 25'd4372, 25'd547, 25'd10712, -25'd11805, -25'd3170, -25'd4263, 25'd9400, -25'd3061}, '{25'd5137, 25'd5247, -25'd10165, -25'd10165, -25'd8526, -25'd3279, 25'd10493, 25'd7214, 25'd5684}, '{25'd3935, -25'd9400, -25'd656, -25'd7870, 25'd5028, 25'd3607, 25'd7433, -25'd4044, 25'd219}, '{25'd2077, -25'd10930, 25'd2186, -25'd11258, -25'd3170, -25'd2077, -25'd4591, -25'd3388, -25'd6777}, '{25'd1312, 25'd6668, -25'd4700, -25'd3498, 25'd5902, 25'd547, -25'd7651, -25'd1530, -25'd8854}, '{-25'd2951, 25'd5465, -25'd10821, 25'd11368, 25'd9619, -25'd3607, -25'd4044, -25'd4154, 25'd7214}, '{25'd7433, 25'd9728, 25'd9072, -25'd8198, -25'd8526, -25'd10930, -25'd4919, 25'd2514, -25'd11586}, '{25'd437, -25'd11586, -25'd4044, -25'd1421, 25'd7433, -25'd5247, -25'd2186, -25'd11040, -25'd5684}, '{25'd2405, -25'd3170, -25'd11805, 25'd1967, -25'd5247, 25'd10603, 25'd2405, -25'd9947, 25'd1967}}, '{'{25'd5465, -25'd2295, 25'd3826, -25'd7542, 25'd11914, -25'd984, 25'd11805, -25'd7323, -25'd109}, '{-25'd6121, 25'd2623, -25'd9619, 25'd13882, 25'd4809, -25'd8635, 25'd1312, 25'd1749, 25'd12789}, '{25'd10930, -25'd6230, 25'd547, -25'd7433, -25'd8744, -25'd5356, 25'd9837, 25'd5356, 25'd2186}, '{25'd11586, -25'd8744, 25'd1967, -25'd9728, 25'd1858, -25'd10056, 25'd3716, -25'd9619, 25'd1749}, '{25'd9072, -25'd5247, -25'd9182, 25'd1749, 25'd2186, 25'd6886, 25'd13117, 25'd11149, -25'd3716}, '{-25'd1749, -25'd1312, 25'd5247, 25'd3716, -25'd4591, 25'd984, -25'd10165, 25'd5793, -25'd3279}, '{-25'd8416, 25'd874, 25'd5137, -25'd6449, 25'd9400, 25'd3279, -25'd6995, 25'd4700, -25'd8198}, '{25'd10493, 25'd6668, 25'd1093, -25'd6995, 25'd3388, -25'd5465, 25'd3498, 25'd6995, -25'd7542}, '{25'd4809, 25'd7323, 25'd1421, 25'd7870, -25'd8963, 25'd12679, -25'd5247, 25'd6230, -25'd6449}}},
    '{'{'{-25'd12327, -25'd4931, -25'd9111, 25'd4824, 25'd5788, 25'd9647, -25'd107, -25'd1501, -25'd10934}, '{-25'd1822, 25'd965, 25'd4073, 25'd7825, 25'd3001, -25'd1822, -25'd9862, 25'd2144, -25'd8468}, '{25'd6432, 25'd4931, 25'd4073, 25'd1286, 25'd3537, -25'd3645, 25'd2894, -25'd2144, -25'd5896}, '{25'd2465, -25'd12863, -25'd10719, 25'd10183, 25'd7503, 25'd9326, -25'd10505, 25'd107, -25'd6110}, '{25'd5360, 25'd536, -25'd8254, 25'd4824, -25'd6646, -25'd10183, -25'd4931, 25'd9433, -25'd4931}, '{25'd2358, 25'd643, -25'd9755, -25'd6860, 25'd2894, -25'd6646, 25'd322, -25'd9755, -25'd9004}, '{25'd2144, -25'd750, -25'd2251, 25'd4395, -25'd4502, 25'd214, -25'd2680, 25'd107, -25'd5360}, '{-25'd8361, 25'd11041, 25'd9219, -25'd8468, 25'd1715, 25'd11684, -25'd2251, -25'd1072, 25'd10934}, '{-25'd5467, -25'd3966, -25'd5145, -25'd8897, 25'd2894, 25'd11148, 25'd0, -25'd4716, -25'd3645}}, '{'{25'd11362, 25'd6324, -25'd4288, 25'd3109, -25'd9755, -25'd6646, -25'd4824, -25'd6003, -25'd6539}, '{25'd13613, -25'd6539, 25'd7932, 25'd2573, 25'd8254, 25'd6003, -25'd9540, 25'd1715, 25'd6432}, '{-25'd6217, -25'd10291, -25'd6432, 25'd1179, 25'd10183, -25'd3859, 25'd5574, -25'd643, 25'd12327}, '{25'd6217, 25'd9540, 25'd7396, -25'd4716, -25'd3216, -25'd6217, -25'd4181, 25'd3109, 25'd7932}, '{-25'd1286, -25'd5788, 25'd10505, -25'd10183, -25'd8039, 25'd10398, 25'd3645, 25'd5681, -25'd7075}, '{25'd429, 25'd6860, -25'd8575, 25'd2573, 25'd3001, 25'd12113, 25'd4395, -25'd7825, 25'd11470}, '{25'd12006, 25'd12756, 25'd6217, -25'd1822, 25'd322, 25'd10398, 25'd10398, -25'd2358, 25'd10505}, '{25'd2358, -25'd10076, 25'd12542, 25'd5896, -25'd9540, 25'd1822, 25'd5467, 25'd11577, 25'd1179}, '{-25'd5896, 25'd12220, 25'd13185, -25'd9969, -25'd7289, -25'd8361, 25'd7825, 25'd10826, -25'd7718}}, '{'{-25'd3109, 25'd1929, 25'd9111, 25'd8468, 25'd11255, 25'd8790, 25'd11362, -25'd10612, 25'd8897}, '{25'd6217, -25'd4181, 25'd1394, 25'd858, -25'd2573, -25'd6432, 25'd8790, -25'd214, -25'd9540}, '{-25'd3430, 25'd5574, -25'd10934, 25'd8897, 25'd5252, -25'd4502, 25'd2251, -25'd3645, 25'd4181}, '{-25'd7289, 25'd2251, 25'd2680, 25'd9004, 25'd429, 25'd536, -25'd7396, 25'd10934, 25'd214}, '{25'd8361, 25'd6539, 25'd1822, -25'd429, 25'd0, -25'd9219, 25'd858, -25'd9111, 25'd9326}, '{25'd3645, 25'd12434, 25'd10719, -25'd8575, -25'd3537, 25'd3216, -25'd2680, 25'd7611, 25'd536}, '{-25'd3109, -25'd8147, 25'd9755, -25'd1715, 25'd11148, -25'd6432, -25'd10612, 25'd10398, 25'd2251}, '{-25'd643, -25'd4716, 25'd3216, -25'd11041, -25'd5896, -25'd5896, 25'd1179, 25'd5681, 25'd5252}, '{-25'd3323, -25'd10398, -25'd3859, -25'd4502, -25'd4824, 25'd4181, -25'd858, -25'd7718, -25'd5681}}},
    '{'{'{25'd5056, 25'd2748, -25'd1209, 25'd10443, 25'd5716, -25'd10663, 25'd3627, -25'd2418, 25'd6595}, '{25'd6485, 25'd10773, -25'd1209, 25'd879, -25'd3737, 25'd2198, -25'd6925, -25'd2198, -25'd5716}, '{25'd2089, 25'd7805, -25'd1869, -25'd6266, 25'd2748, 25'd5606, -25'd6815, -25'd1319, 25'd10773}, '{25'd10882, 25'd3737, 25'd8244, -25'd5056, -25'd1869, -25'd6815, 25'd7805, 25'd4287, -25'd7145}, '{-25'd2638, -25'd7695, -25'd11432, -25'd9014, 25'd1869, 25'd7805, 25'd8024, -25'd2089, -25'd6815}, '{25'd6376, -25'd11432, -25'd9124, -25'd769, 25'd11652, 25'd11872, -25'd10553, -25'd2748, -25'd6705}, '{-25'd1429, 25'd1429, 25'd6595, -25'd8684, 25'd10992, 25'd9783, -25'd989, 25'd10003, 25'd9014}, '{25'd2528, -25'd8244, 25'd3737, 25'd10223, 25'd9124, 25'd7475, 25'd7365, -25'd1319, -25'd9124}, '{25'd5276, -25'd5056, -25'd2198, 25'd660, 25'd3627, 25'd3188, 25'd4837, -25'd220, 25'd3518}}, '{'{25'd11322, -25'd1649, -25'd3737, 25'd2308, -25'd8574, 25'd330, -25'd5276, 25'd9893, 25'd10992}, '{25'd11872, -25'd1649, 25'd10443, 25'd4067, 25'd4397, -25'd4617, 25'd7365, -25'd7695, -25'd11212}, '{25'd11542, 25'd6485, -25'd660, -25'd7805, 25'd330, 25'd1209, -25'd5166, 25'd9893, -25'd10333}, '{25'd3078, -25'd1649, -25'd8134, 25'd9234, 25'd6595, 25'd1649, -25'd4617, 25'd2748, 25'd220}, '{25'd6156, 25'd7805, -25'd5166, 25'd13960, 25'd110, 25'd6485, 25'd8794, -25'd4287, 25'd11102}, '{25'd7475, -25'd7805, -25'd6485, -25'd10773, -25'd660, -25'd4507, -25'd11872, -25'd3957, -25'd7035}, '{25'd2858, -25'd8464, -25'd1539, 25'd4837, 25'd10333, -25'd5276, 25'd7915, -25'd8244, 25'd8464}, '{-25'd4507, -25'd5936, 25'd10553, -25'd1539, 25'd11762, -25'd4287, -25'd1979, -25'd3847, -25'd5936}, '{-25'd5276, -25'd2198, -25'd2198, -25'd220, -25'd4947, -25'd10663, -25'd11432, -25'd1209, -25'd1759}}, '{'{25'd1759, 25'd5826, -25'd9893, 25'd769, 25'd10992, -25'd5276, 25'd10663, -25'd440, 25'd550}, '{-25'd7035, 25'd12092, 25'd6485, -25'd1979, 25'd10223, 25'd11102, -25'd5496, 25'd5826, 25'd12641}, '{-25'd7475, 25'd10553, -25'd5826, 25'd5166, -25'd5936, -25'd5056, -25'd8794, 25'd6266, 25'd9453}, '{-25'd5826, 25'd3847, -25'd2748, 25'd9234, 25'd7475, 25'd8354, 25'd5056, 25'd11652, -25'd4727}, '{25'd9893, 25'd4837, -25'd3078, -25'd6705, -25'd7805, -25'd4397, -25'd4507, -25'd5386, -25'd3518}, '{25'd4727, 25'd440, -25'd2638, 25'd1979, 25'd10223, -25'd3078, -25'd4727, 25'd2748, -25'd3737}, '{25'd2748, 25'd4177, 25'd4177, -25'd6376, -25'd7365, 25'd1869, -25'd8134, -25'd5826, -25'd5496}, '{-25'd4397, -25'd7475, 25'd10773, 25'd7585, 25'd0, -25'd1539, 25'd11982, -25'd4397, 25'd879}, '{-25'd879, 25'd12311, -25'd9014, 25'd2968, 25'd12861, 25'd6705, -25'd9893, -25'd2968, -25'd8794}}},
    '{'{'{25'd9035, 25'd9263, 25'd4231, -25'd1258, -25'd11550, -25'd10979, 25'd10178, -25'd3545, -25'd8120}, '{-25'd5832, 25'd3316, -25'd9606, -25'd1601, 25'd7891, 25'd5261, -25'd5375, -25'd6519, -25'd1830}, '{-25'd1029, 25'd5146, 25'd1029, 25'd11550, -25'd3888, -25'd2287, 25'd6633, -25'd3888, 25'd4918}, '{-25'd686, -25'd4117, 25'd11665, -25'd1487, 25'd6976, -25'd3431, -25'd7090, -25'd1029, -25'd10292}, '{-25'd9949, 25'd3202, -25'd2058, 25'd9949, 25'd2516, -25'd229, 25'd11436, 25'd12351, -25'd4460}, '{25'd1944, -25'd7090, -25'd11436, -25'd4689, 25'd6862, -25'd6061, -25'd915, -25'd4460, 25'd7891}, '{-25'd10750, -25'd8577, 25'd10864, 25'd801, -25'd5489, -25'd3888, -25'd9263, 25'd8120, -25'd9949}, '{-25'd11207, 25'd10178, -25'd6061, 25'd2058, -25'd5718, -25'd7090, -25'd7548, -25'd8691, 25'd915}, '{-25'd1830, -25'd3545, -25'd3088, -25'd10407, -25'd10521, 25'd3545, -25'd2973, -25'd114, -25'd3316}}, '{'{-25'd915, -25'd13495, -25'd3888, 25'd3088, -25'd7548, 25'd457, -25'd229, 25'd1944, 25'd4003}, '{-25'd229, -25'd4117, -25'd10064, -25'd13495, -25'd7777, 25'd4918, -25'd9492, -25'd12237, 25'd9035}, '{-25'd14409, 25'd4803, 25'd7319, -25'd13723, -25'd2516, 25'd2173, -25'd5032, -25'd12465, 25'd8120}, '{-25'd6519, 25'd7433, 25'd8577, 25'd8348, -25'd9835, -25'd6061, 25'd8463, -25'd8691, -25'd4574}, '{25'd4346, 25'd6175, -25'd4346, -25'd4574, 25'd4689, 25'd8348, -25'd10636, 25'd8120, -25'd12694}, '{25'd8920, 25'd5718, 25'd114, -25'd10979, -25'd12580, -25'd11550, -25'd10864, -25'd11207, -25'd1372}, '{-25'd13838, -25'd7205, -25'd8348, -25'd1144, -25'd6290, 25'd6519, -25'd114, -25'd5604, -25'd2630}, '{25'd5832, 25'd2859, -25'd13266, 25'd6633, -25'd11779, -25'd9378, 25'd3545, 25'd2745, -25'd6862}, '{25'd4803, -25'd457, -25'd9492, 25'd572, -25'd7662, -25'd5947, -25'd801, -25'd10292, -25'd5832}}, '{'{25'd6747, 25'd114, -25'd7205, -25'd3545, 25'd6061, 25'd6404, 25'd10979, 25'd0, 25'd1487}, '{25'd10407, -25'd1029, 25'd6747, -25'd1487, -25'd6519, -25'd4689, 25'd14524, 25'd5832, -25'd6747}, '{-25'd3774, 25'd13151, 25'd12008, 25'd915, 25'd5604, 25'd14066, 25'd12008, 25'd4574, -25'd5146}, '{-25'd5718, 25'd5947, -25'd6633, 25'd0, 25'd229, 25'd343, 25'd5146, 25'd7205, 25'd8234}, '{25'd12008, -25'd915, 25'd5832, 25'd1944, 25'd1715, 25'd13723, -25'd8120, -25'd5032, 25'd12122}, '{25'd1715, -25'd2058, -25'd8005, 25'd8463, 25'd13266, 25'd9721, -25'd5832, -25'd2287, 25'd7205}, '{25'd11550, 25'd11779, 25'd3888, -25'd4346, 25'd6061, 25'd12237, 25'd8120, 25'd801, 25'd2516}, '{25'd7777, 25'd4460, 25'd5489, 25'd915, 25'd11779, 25'd11779, 25'd13838, 25'd5146, -25'd3774}, '{25'd5375, 25'd343, -25'd1487, 25'd11322, 25'd9606, -25'd6404, -25'd7090, 25'd14409, 25'd2287}}},
    '{'{'{-25'd4826, -25'd4203, 25'd3269, -25'd1557, 25'd11208, 25'd6382, -25'd5604, 25'd2491, 25'd6227}, '{-25'd1868, 25'd3892, 25'd3892, 25'd10741, -25'd2024, 25'd1712, -25'd7472, -25'd8717, -25'd4670}, '{-25'd10741, 25'd10430, 25'd6227, -25'd2802, 25'd7316, -25'd7472, 25'd12142, -25'd3425, 25'd10118}, '{25'd10274, -25'd11052, -25'd3736, 25'd9340, 25'd3269, 25'd11364, 25'd3269, 25'd5760, 25'd8250}, '{25'd10897, 25'd3736, 25'd10118, 25'd10741, -25'd3892, -25'd8873, 25'd11831, -25'd7005, -25'd5604}, '{25'd934, 25'd7628, 25'd14633, -25'd7783, -25'd2646, -25'd6538, -25'd4359, -25'd6694, 25'd8095}, '{25'd10741, -25'd8873, 25'd1868, -25'd467, -25'd2024, -25'd311, 25'd11208, -25'd1712, 25'd8406}, '{25'd6071, 25'd3892, -25'd7161, -25'd3113, -25'd2491, -25'd8095, 25'd1868, 25'd11986, 25'd4514}, '{25'd311, 25'd6538, -25'd1712, -25'd7472, -25'd6382, -25'd5915, 25'd9807, -25'd7472, -25'd6382}}, '{'{-25'd9340, -25'd11831, -25'd10430, -25'd10897, -25'd15722, -25'd4359, 25'd2646, 25'd5760, -25'd14166}, '{-25'd19769, 25'd311, 25'd4047, 25'd5137, -25'd13543, 25'd1090, -25'd12298, -25'd5137, -25'd8562}, '{-25'd1245, -25'd3113, 25'd4203, -25'd2646, -25'd13387, -25'd15878, -25'd1090, -25'd9963, 25'd5293}, '{-25'd2335, -25'd14944, -25'd7783, -25'd14944, -25'd11364, -25'd1712, -25'd3269, -25'd8250, -25'd9029}, '{-25'd5137, -25'd13543, -25'd15722, -25'd16033, -25'd12920, 25'd2958, -25'd14633, -25'd16345, -25'd2646}, '{25'd5915, -25'd12920, -25'd2335, -25'd2491, -25'd10897, -25'd5448, 25'd5137, -25'd12298, 25'd2958}, '{-25'd14788, 25'd1401, 25'd6694, -25'd2179, -25'd10430, -25'd5604, -25'd1868, -25'd14477, -25'd1090}, '{-25'd14166, -25'd5760, -25'd13232, 25'd4981, -25'd8562, 25'd4826, -25'd12142, -25'd778, -25'd12920}, '{-25'd6227, -25'd12765, -25'd11052, 25'd467, 25'd3269, -25'd4047, 25'd9029, -25'd10741, -25'd10118}}, '{'{25'd7316, 25'd1245, 25'd8717, -25'd5137, 25'd11831, 25'd11986, 25'd7472, 25'd7783, 25'd2646}, '{25'd6227, 25'd2179, 25'd1557, 25'd8717, 25'd5915, 25'd6694, 25'd12142, -25'd6071, 25'd14166}, '{25'd2958, 25'd13543, -25'd3892, 25'd9029, 25'd4203, 25'd16189, -25'd2491, 25'd14477, 25'd8095}, '{-25'd3113, 25'd5137, -25'd6538, 25'd156, -25'd467, 25'd7783, -25'd3113, -25'd934, 25'd2491}, '{-25'd2958, 25'd156, -25'd156, -25'd4203, -25'd934, 25'd11831, 25'd1401, -25'd1868, 25'd16033}, '{25'd10118, -25'd467, 25'd4359, -25'd1868, 25'd16656, 25'd3113, -25'd4359, 25'd3892, 25'd10274}, '{25'd14010, 25'd8562, 25'd7628, -25'd2335, 25'd9496, 25'd2958, 25'd311, -25'd4359, 25'd11519}, '{25'd10274, 25'd11675, 25'd15099, 25'd16345, 25'd2335, 25'd3892, -25'd5293, -25'd1245, 25'd11208}, '{-25'd5915, 25'd6071, 25'd1401, 25'd4203, -25'd623, -25'd1245, -25'd467, -25'd1401, 25'd13854}}},
    '{'{'{25'd8653, 25'd5421, 25'd2398, 25'd5421, 25'd3023, 25'd521, -25'd938, -25'd1564, -25'd1460}, '{25'd12615, -25'd10634, -25'd5943, 25'd12615, 25'd626, -25'd2398, -25'd8653, 25'd1668, -25'd10530}, '{-25'd4379, -25'd417, 25'd2711, -25'd2398, -25'd1668, -25'd4587, 25'd521, -25'd4587, 25'd10634}, '{-25'd2711, -25'd11155, 25'd6151, -25'd6568, 25'd5109, 25'd2502, -25'd3023, 25'd7923, 25'd5213}, '{25'd6881, 25'd10843, 25'd8445, 25'd2606, 25'd6985, -25'd9800, 25'd11364, 25'd4900, 25'd1877}, '{25'd4900, -25'd2189, -25'd8653, 25'd3649, 25'd2502, -25'd3857, 25'd104, 25'd209, -25'd1460}, '{-25'd9487, 25'd6151, -25'd3753, 25'd2294, 25'd3128, -25'd8132, -25'd1043, -25'd5734, -25'd3232}, '{-25'd9904, -25'd1981, 25'd10738, 25'd2919, -25'd8445, 25'd4900, 25'd4900, 25'd2085, -25'd3753}, '{-25'd6985, -25'd5734, -25'd5004, 25'd3232, -25'd6151, -25'd9279, -25'd12094, -25'd8757, -25'd11260}}, '{'{25'd6881, 25'd9383, -25'd13032, 25'd4066, 25'd5734, -25'd4170, -25'd834, -25'd10426, 25'd2711}, '{25'd1564, -25'd6881, -25'd8757, -25'd6672, 25'd6360, -25'd11781, -25'd9487, -25'd11260, -25'd209}, '{25'd8549, 25'd9904, -25'd730, 25'd8340, -25'd8966, -25'd1668, 25'd5630, -25'd209, -25'd1877}, '{25'd9279, 25'd9279, 25'd10947, 25'd5526, -25'd730, 25'd2815, -25'd12302, 25'd104, 25'd2398}, '{-25'd5526, -25'd3440, -25'd10530, 25'd5213, -25'd5317, 25'd0, -25'd5943, 25'd10634, 25'd209}, '{-25'd8340, -25'd12615, 25'd8340, 25'd11260, 25'd6151, 25'd10738, 25'd7611, 25'd9800, -25'd1668}, '{25'd6464, -25'd8653, 25'd10530, 25'd10738, -25'd11155, -25'd12928, -25'd5317, -25'd6047, -25'd6985}, '{-25'd12198, -25'd2294, -25'd7923, -25'd8445, -25'd6777, 25'd5317, -25'd4691, -25'd4691, -25'd3336}, '{-25'd1251, 25'd9591, -25'd7715, -25'd3962, 25'd1043, -25'd4587, -25'd9279, 25'd10008, -25'd6047}}, '{'{25'd834, -25'd9279, -25'd6568, -25'd1355, 25'd8549, 25'd5734, 25'd6672, 25'd626, 25'd6047}, '{25'd6464, -25'd2189, -25'd7819, -25'd1668, 25'd7611, 25'd626, -25'd3023, 25'd313, 25'd2815}, '{-25'd7194, -25'd2711, 25'd8549, -25'd5526, -25'd8132, -25'd3962, 25'd2606, -25'd1772, -25'd7611}, '{-25'd1043, -25'd1564, 25'd11364, 25'd1981, -25'd7819, -25'd4379, -25'd9696, -25'd9383, -25'd8236}, '{-25'd3962, -25'd11364, 25'd9070, -25'd8132, -25'd6672, 25'd2085, 25'd4170, 25'd8028, 25'd2189}, '{-25'd4483, -25'd11364, 25'd6360, 25'd7402, -25'd3336, -25'd8757, -25'd8028, 25'd10738, -25'd6985}, '{-25'd4066, 25'd10321, 25'd10008, -25'd4900, 25'd10321, -25'd6360, 25'd6464, 25'd1981, -25'd4587}, '{25'd5734, -25'd10947, -25'd9383, -25'd7715, 25'd11051, -25'd11468, 25'd10217, 25'd12719, 25'd13240}, '{25'd4379, 25'd1147, 25'd2085, 25'd9800, -25'd4691, 25'd11051, 25'd10634, -25'd3649, 25'd8757}}},
    '{'{'{25'd8097, 25'd3216, 25'd1331, -25'd887, -25'd3882, 25'd3771, -25'd8540, 25'd2329, 25'd0}, '{-25'd1775, -25'd4991, 25'd555, 25'd3327, 25'd5656, 25'd4215, 25'd10426, 25'd10648, -25'd3882}, '{25'd4769, 25'd5213, -25'd9538, -25'd3549, 25'd5656, 25'd222, -25'd9871, -25'd1442, -25'd7542}, '{-25'd11313, -25'd998, 25'd9982, 25'd9206, -25'd3549, 25'd111, 25'd10426, -25'd4215, -25'd6433}, '{-25'd5656, 25'd6877, -25'd4547, -25'd1996, -25'd4769, 25'd2329, 25'd10648, -25'd7431, 25'd2662}, '{-25'd6433, 25'd9538, -25'd5767, 25'd3993, 25'd5546, 25'd776, -25'd2551, 25'd5102, 25'd2551}, '{-25'd4547, 25'd3549, -25'd6100, 25'd4326, 25'd8873, -25'd7986, 25'd10426, -25'd11424, -25'd1664}, '{-25'd5324, 25'd11091, -25'd10315, 25'd1553, -25'd10204, -25'd10980, 25'd444, -25'd9649, -25'd7653}, '{25'd8097, 25'd3993, -25'd10537, -25'd8429, -25'd11202, 25'd11313, -25'd2551, -25'd3660, -25'd222}}, '{'{25'd14086, -25'd1553, -25'd6877, 25'd4326, 25'd12200, -25'd9982, -25'd2662, 25'd1331, 25'd12089}, '{25'd111, 25'd10758, -25'd8540, -25'd6655, 25'd3216, 25'd998, -25'd5546, 25'd4991, -25'd3327}, '{25'd4880, -25'd2551, 25'd4436, 25'd555, 25'd11424, 25'd10426, 25'd6544, 25'd3106, -25'd6766}, '{25'd776, -25'd4991, -25'd4658, -25'd5102, 25'd10869, -25'd7986, -25'd2440, -25'd10869, 25'd5767}, '{25'd9538, 25'd5989, 25'd5435, 25'd1775, -25'd8984, 25'd1885, -25'd1996, -25'd8318, -25'd7209}, '{25'd5213, -25'd1109, 25'd4547, 25'd10648, 25'd9538, -25'd6987, 25'd7320, 25'd0, 25'd11424}, '{25'd1775, 25'd11202, 25'd13198, -25'd2218, 25'd11646, 25'd7098, 25'd4769, -25'd5989, -25'd2773}, '{25'd10537, 25'd11424, -25'd6211, -25'd4104, 25'd5213, -25'd555, -25'd10093, -25'd10537, -25'd11091}, '{25'd10648, -25'd5324, 25'd333, 25'd9427, 25'd7320, 25'd665, 25'd8207, 25'd4547, -25'd10758}}, '{'{-25'd8984, -25'd998, 25'd7209, 25'd555, 25'd6766, -25'd2218, -25'd2218, -25'd2884, -25'd6322}, '{-25'd776, -25'd11535, 25'd2107, 25'd1220, 25'd8097, -25'd555, 25'd222, 25'd2995, -25'd5767}, '{-25'd8207, -25'd1553, -25'd6100, -25'd6655, 25'd4658, -25'd11646, 25'd5324, 25'd3993, -25'd6544}, '{-25'd3327, -25'd776, 25'd7209, -25'd1442, 25'd5767, 25'd7875, -25'd998, 25'd5989, 25'd4104}, '{-25'd1331, 25'd3327, 25'd8873, 25'd10204, 25'd2551, -25'd1331, 25'd3438, 25'd7431, -25'd11091}, '{-25'd8429, -25'd444, -25'd2551, 25'd1220, -25'd4326, 25'd8984, 25'd333, 25'd1775, 25'd8318}, '{-25'd2218, 25'd3882, -25'd4326, -25'd6322, -25'd6766, 25'd7542, -25'd8429, 25'd5878, -25'd10758}, '{-25'd1553, 25'd4880, -25'd6766, 25'd12755, -25'd1109, -25'd8318, -25'd5656, 25'd2551, 25'd4215}, '{25'd9317, 25'd11313, -25'd2995, 25'd8873, 25'd3993, -25'd8984, -25'd5767, 25'd7209, -25'd3993}}},
    '{'{'{-25'd8607, 25'd4616, 25'd4241, -25'd8483, -25'd3243, 25'd7111, 25'd624, 25'd8483, -25'd10728}, '{25'd9980, -25'd4616, 25'd3992, -25'd10603, -25'd4616, -25'd10229, 25'd3618, -25'd9231, 25'd10479}, '{25'd9855, -25'd3368, 25'd1123, 25'd8857, -25'd2994, -25'd8607, 25'd12475, 25'd12475, 25'd0}, '{25'd5239, -25'd10229, 25'd10104, 25'd3992, 25'd1372, 25'd2121, -25'd3992, -25'd4117, 25'd4865}, '{25'd3493, 25'd10354, -25'd4366, 25'd11227, 25'd1746, 25'd4241, 25'd0, -25'd10479, 25'd7485}, '{-25'd374, -25'd8483, -25'd5115, 25'd12100, -25'd5115, -25'd1871, -25'd7111, -25'd2869, 25'd2495}, '{25'd10229, -25'd7610, 25'd3243, -25'd10479, -25'd998, -25'd8233, -25'd6612, 25'd5863, -25'd7360}, '{25'd2620, 25'd11976, 25'd1247, -25'd9730, 25'd1622, 25'd4740, -25'd7859, -25'd9106, -25'd7610}, '{-25'd6861, 25'd5115, -25'd1871, 25'd9481, 25'd12974, -25'd5115, -25'd3368, -25'd3992, 25'd7859}}, '{'{-25'd5115, 25'd10853, 25'd1123, -25'd5239, 25'd8358, 25'd8483, 25'd15843, 25'd11227, -25'd249}, '{25'd7485, -25'd4616, -25'd7235, 25'd9231, 25'd7610, -25'd2994, 25'd4117, 25'd9481, 25'd15593}, '{25'd2994, 25'd1123, 25'd8483, -25'd7360, 25'd7859, 25'd12350, 25'd15843, 25'd11851, 25'd2245}, '{25'd125, -25'd873, 25'd9106, 25'd13348, -25'd4241, 25'd13722, 25'd9855, 25'd10104, 25'd13223}, '{25'd4491, -25'd1622, 25'd8483, -25'd5489, 25'd1996, 25'd12849, 25'd11477, 25'd1123, -25'd2121}, '{25'd12225, -25'd2620, 25'd3119, 25'd4241, 25'd2370, 25'd6861, 25'd11227, -25'd7859, -25'd8109}, '{25'd5115, -25'd125, -25'd5489, -25'd1622, 25'd873, -25'd998, 25'd7360, 25'd2121, 25'd11726}, '{-25'd125, -25'd4491, -25'd8483, 25'd3742, 25'd9980, -25'd5115, -25'd8109, -25'd8607, 25'd14221}, '{25'd12974, -25'd9106, 25'd4865, -25'd9605, 25'd4740, 25'd624, 25'd12849, 25'd5988, 25'd2994}}, '{'{-25'd3867, 25'd3618, 25'd6861, -25'd5364, 25'd873, 25'd1871, 25'd6113, -25'd9855, -25'd11601}, '{-25'd3493, -25'd7984, -25'd4117, 25'd3493, 25'd8857, 25'd6113, 25'd6113, -25'd8607, -25'd2744}, '{25'd3742, -25'd2495, -25'd8732, -25'd5489, -25'd7235, 25'd6237, 25'd8982, 25'd3742, -25'd4616}, '{-25'd1746, -25'd7610, -25'd7610, -25'd2994, -25'd4117, 25'd8732, -25'd7859, -25'd9231, 25'd7610}, '{-25'd6113, 25'd1996, -25'd3368, -25'd11102, -25'd1622, -25'd4740, -25'd11227, 25'd6237, -25'd4616}, '{-25'd4616, 25'd9855, -25'd873, 25'd125, 25'd4117, 25'd8982, -25'd1996, -25'd11477, 25'd6487}, '{25'd6237, -25'd5364, -25'd2620, 25'd12350, 25'd4117, 25'd2245, -25'd9106, 25'd3992, 25'd8607}, '{-25'd7360, -25'd8732, -25'd7360, 25'd4366, -25'd8982, 25'd2370, 25'd7485, 25'd3618, 25'd6113}, '{-25'd5988, 25'd1372, 25'd748, -25'd6986, -25'd6487, 25'd2620, 25'd873, -25'd6986, 25'd0}}},
    '{'{'{25'd10033, 25'd6337, 25'd8660, 25'd9822, -25'd3063, -25'd6125, -25'd10456, 25'd422, 25'd4964}, '{25'd4753, -25'd2112, 25'd5597, -25'd3696, 25'd12145, 25'd4858, -25'd6231, -25'd2218, 25'd6654}, '{-25'd9188, 25'd6125, -25'd9294, 25'd2323, -25'd7182, 25'd6337, 25'd634, -25'd9928, -25'd8343}, '{-25'd6442, -25'd3274, 25'd951, 25'd7287, -25'd4013, -25'd8977, 25'd10667, 25'd9188, -25'd3591}, '{25'd2852, -25'd3063, 25'd7710, -25'd1795, -25'd9188, 25'd7815, -25'd845, -25'd6020, -25'd211}, '{25'd9399, 25'd1479, 25'd3696, 25'd9083, -25'd6337, -25'd317, 25'd8238, -25'd3696, 25'd7921}, '{25'd11406, -25'd2007, 25'd6548, 25'd7287, -25'd3908, 25'd8343, 25'd9611, -25'd8343, -25'd5914}, '{25'd2218, -25'd4753, -25'd8027, -25'd1795, -25'd4436, -25'd2746, 25'd3696, 25'd1373, 25'd10139}, '{25'd6759, -25'd9928, 25'd317, 25'd4330, 25'd8132, -25'd9822, -25'd11300, -25'd3591, 25'd9188}}, '{'{-25'd6865, 25'd2112, -25'd6020, 25'd8977, 25'd6865, 25'd8449, -25'd5809, -25'd1795, 25'd3274}, '{-25'd11934, -25'd7815, -25'd8449, 25'd2007, 25'd7287, 25'd9928, 25'd8555, -25'd9928, -25'd3274}, '{-25'd8871, -25'd10244, -25'd7393, -25'd12673, -25'd4330, 25'd6654, 25'd8343, 25'd3380, 25'd3802}, '{25'd6231, -25'd528, 25'd5175, 25'd0, -25'd4858, 25'd0, -25'd4119, -25'd106, -25'd9188}, '{-25'd3485, 25'd6970, -25'd8343, 25'd6125, 25'd8449, -25'd845, -25'd7710, 25'd739, 25'd951}, '{-25'd9505, 25'd7076, -25'd12885, -25'd13413, 25'd7815, 25'd2007, 25'd5809, 25'd8238, 25'd5492}, '{-25'd11617, 25'd6970, 25'd6759, 25'd9716, 25'd9611, -25'd11089, 25'd422, -25'd6020, -25'd2007}, '{25'd1795, -25'd10878, 25'd3168, 25'd6548, -25'd8555, -25'd11512, 25'd951, -25'd10667, 25'd2640}, '{25'd634, -25'd7393, 25'd4119, -25'd7815, 25'd5597, -25'd739, -25'd739, -25'd528, 25'd6865}}, '{'{25'd6654, 25'd5281, 25'd2852, -25'd3591, -25'd5281, -25'd3485, 25'd12885, -25'd106, -25'd8871}, '{-25'd4858, 25'd12779, -25'd5386, 25'd6865, 25'd3485, -25'd8027, 25'd1584, 25'd9822, -25'd9611}, '{25'd2429, -25'd10456, -25'd2535, 25'd8449, -25'd5281, -25'd5386, 25'd10244, 25'd3908, -25'd7815}, '{25'd9399, 25'd4753, 25'd4858, 25'd1690, 25'd12251, 25'd11617, 25'd7815, 25'd2429, 25'd8871}, '{-25'd2957, -25'd8766, 25'd12251, 25'd2957, 25'd9083, 25'd1795, 25'd8238, -25'd6020, 25'd11406}, '{25'd1479, -25'd317, -25'd1479, -25'd1267, 25'd8132, -25'd528, 25'd1479, -25'd3380, 25'd2746}, '{25'd5386, -25'd1901, 25'd11512, -25'd10139, 25'd4541, 25'd9505, 25'd10456, -25'd7815, 25'd5386}, '{-25'd1584, 25'd739, 25'd1162, 25'd5069, 25'd11934, 25'd3696, -25'd3591, 25'd9611, 25'd7498}, '{-25'd8238, 25'd9716, 25'd8766, 25'd8766, 25'd10139, 25'd10667, -25'd10139, -25'd2746, 25'd11617}}},
    '{'{'{-25'd5118, -25'd7949, 25'd8058, -25'd1742, 25'd218, 25'd10562, 25'd5771, 25'd5227, 25'd10454}, '{25'd1851, 25'd5771, 25'd4900, 25'd762, -25'd4356, 25'd7513, -25'd327, 25'd1960, -25'd5336}, '{25'd5989, -25'd1742, 25'd871, 25'd7731, 25'd0, -25'd11216, 25'd8167, 25'd3158, -25'd3376}, '{-25'd9038, -25'd4682, -25'd7405, -25'd6316, 25'd2722, -25'd1307, 25'd436, -25'd10018, 25'd4682}, '{-25'd2178, -25'd2722, 25'd9691, 25'd6098, 25'd8820, 25'd8058, 25'd6642, 25'd9365, -25'd8385}, '{-25'd109, -25'd7296, 25'd10018, 25'd1416, -25'd4900, -25'd2722, 25'd9909, 25'd7622, -25'd4138}, '{-25'd5445, 25'd11760, 25'd218, 25'd327, 25'd980, 25'd6207, -25'd5771, 25'd1524, -25'd1198}, '{25'd1633, 25'd8058, -25'd2069, 25'd8602, 25'd1416, -25'd9147, 25'd980, -25'd11760, -25'd1307}, '{-25'd5009, -25'd1960, -25'd2831, 25'd8058, -25'd3593, -25'd9365, -25'd7622, -25'd10345, -25'd9582}}, '{'{-25'd5445, -25'd6425, -25'd1416, 25'd5336, 25'd109, -25'd10345, -25'd7840, 25'd1089, -25'd3811}, '{-25'd6969, 25'd9691, 25'd1633, -25'd544, -25'd4465, -25'd10889, -25'd327, 25'd4900, 25'd2287}, '{25'd10562, 25'd1742, 25'd7187, 25'd5989, -25'd5009, -25'd6316, 25'd2178, 25'd5445, 25'd9038}, '{-25'd8929, 25'd9365, 25'd8711, -25'd7187, -25'd3811, -25'd3811, -25'd10671, 25'd2613, -25'd2287}, '{-25'd3485, -25'd8385, 25'd11760, 25'd4465, 25'd1851, 25'd980, 25'd9909, 25'd7513, -25'd1960}, '{-25'd2069, 25'd1307, 25'd4465, 25'd6533, -25'd8276, 25'd10127, 25'd11869, -25'd9909, 25'd10345}, '{25'd5336, 25'd2178, 25'd11869, 25'd6316, 25'd5662, 25'd5553, 25'd1742, -25'd10889, -25'd9691}, '{25'd6751, -25'd3158, 25'd5336, 25'd12196, -25'd6207, -25'd2613, 25'd1851, 25'd10236, -25'd8167}, '{25'd1633, -25'd8820, -25'd1524, 25'd12196, -25'd4791, 25'd13829, 25'd2178, -25'd11107, 25'd7078}}, '{'{25'd1851, 25'd3702, 25'd5445, -25'd1416, 25'd11542, -25'd7078, 25'd10780, -25'd3049, 25'd1633}, '{25'd2504, 25'd4791, -25'd10780, 25'd5227, -25'd10236, -25'd5989, -25'd9582, 25'd11107, 25'd1742}, '{-25'd4356, -25'd1633, 25'd8058, 25'd1416, -25'd4900, -25'd3049, -25'd4791, -25'd2396, 25'd6860}, '{-25'd6207, 25'd6098, -25'd8820, -25'd1633, -25'd7949, -25'd2069, 25'd7405, -25'd1198, 25'd5009}, '{-25'd218, -25'd5662, -25'd9474, 25'd6642, -25'd109, -25'd2722, -25'd4573, 25'd3920, 25'd8167}, '{25'd6751, -25'd5989, -25'd2504, -25'd5880, 25'd11651, 25'd6207, -25'd3811, -25'd6098, 25'd980}, '{25'd4465, 25'd3049, 25'd7949, 25'd6751, -25'd6969, 25'd980, -25'd1851, -25'd6425, -25'd8711}, '{-25'd6316, 25'd11216, 25'd0, 25'd3267, -25'd653, 25'd9256, -25'd6642, 25'd9365, 25'd9800}, '{-25'd9038, 25'd3267, -25'd3049, 25'd1851, -25'd6751, -25'd8711, 25'd1633, -25'd2940, -25'd1851}}},
    '{'{'{25'd6894, 25'd5709, -25'd2585, 25'd10988, 25'd646, 25'd2585, -25'd2047, 25'd0, 25'd3878}, '{-25'd9588, -25'd7649, 25'd215, 25'd4848, 25'd5279, 25'd9157, -25'd5925, -25'd1400, -25'd108}, '{-25'd2478, -25'd7433, -25'd1185, -25'd7972, -25'd9372, -25'd3124, 25'd11096, -25'd3232, 25'd3770}, '{-25'd11096, -25'd1831, 25'd108, -25'd4524, 25'd11634, -25'd4632, -25'd2155, 25'd11096, -25'd10342}, '{25'd431, 25'd10234, 25'd6571, -25'd1508, 25'd3770, -25'd4201, -25'd9049, 25'd7864, 25'd11742}, '{-25'd6464, -25'd970, -25'd7218, 25'd8941, -25'd7002, -25'd9695, -25'd8510, -25'd7756, 25'd3986}, '{25'd1724, 25'd11311, -25'd6248, 25'd2155, 25'd11096, -25'd8726, -25'd3986, -25'd6248, -25'd6356}, '{25'd9911, 25'd3232, 25'd3878, 25'd7864, -25'd7325, 25'd9480, -25'd11096, 25'd431, -25'd10773}, '{-25'd5709, 25'd11096, 25'd3124, 25'd2262, 25'd8079, 25'd6140, -25'd2693, -25'd6464, 25'd0}}, '{'{25'd6248, 25'd10126, -25'd1831, -25'd646, 25'd2801, 25'd10018, -25'd3555, 25'd4524, -25'd215}, '{-25'd5925, -25'd6787, 25'd1939, 25'd2155, 25'd5602, -25'd9588, 25'd11742, 25'd7433, 25'd8079}, '{-25'd12065, -25'd539, -25'd2155, -25'd3555, -25'd7541, -25'd7649, 25'd1185, -25'd6140, 25'd7864}, '{25'd970, -25'd6140, -25'd11527, -25'd4524, 25'd3986, 25'd10665, 25'd9049, 25'd4417, 25'd6356}, '{-25'd754, -25'd3447, 25'd9803, 25'd11096, 25'd10018, 25'd5494, 25'd9264, -25'd323, -25'd2155}, '{25'd7972, 25'd3447, -25'd8726, 25'd4740, -25'd4201, 25'd1616, -25'd2370, 25'd7433, -25'd2801}, '{25'd10234, -25'd7649, -25'd646, -25'd1508, 25'd1616, 25'd862, 25'd5279, -25'd2909, 25'd11096}, '{-25'd5386, 25'd3878, 25'd1400, -25'd1831, -25'd3124, 25'd1724, -25'd7649, 25'd2478, 25'd4524}, '{-25'd2047, 25'd8726, 25'd9049, 25'd1939, 25'd4094, -25'd9157, 25'd2262, -25'd6140, -25'd10018}}, '{'{-25'd862, 25'd10234, -25'd970, -25'd6894, -25'd7972, 25'd7325, -25'd2801, -25'd3770, -25'd4524}, '{25'd11419, 25'd6033, -25'd4524, -25'd3447, -25'd2801, 25'd7972, 25'd10557, -25'd2585, 25'd11096}, '{-25'd3770, 25'd11958, -25'd970, -25'd4955, 25'd4201, 25'd1293, -25'd7649, 25'd5709, 25'd7110}, '{-25'd754, 25'd4094, -25'd1400, -25'd6140, -25'd6248, -25'd3663, -25'd6787, -25'd1293, 25'd9049}, '{25'd4417, 25'd3339, 25'd4309, -25'd3016, -25'd215, 25'd6894, -25'd2585, 25'd2155, 25'd10449}, '{25'd8079, 25'd215, 25'd1616, 25'd3339, 25'd3663, -25'd6248, 25'd10557, -25'd1616, -25'd9588}, '{25'd7002, 25'd11742, -25'd10773, -25'd6571, -25'd10773, -25'd9049, -25'd9803, -25'd1616, -25'd3770}, '{-25'd4309, -25'd9480, -25'd4740, 25'd10342, -25'd1077, 25'd11850, -25'd9911, 25'd7110, 25'd13681}, '{25'd5279, -25'd9803, 25'd6679, -25'd215, 25'd6033, -25'd3555, -25'd9372, 25'd6464, 25'd6464}}},
    '{'{'{25'd9896, -25'd6597, 25'd11157, -25'd10187, -25'd6694, -25'd7955, 25'd4560, 25'd4560, 25'd8149}, '{25'd2619, 25'd6306, 25'd3105, 25'd5239, -25'd970, 25'd3493, 25'd1746, 25'd2037, 25'd2910}, '{25'd970, -25'd1940, 25'd11545, -25'd5045, -25'd5336, -25'd7373, -25'd6985, 25'd5045, 25'd11060}, '{25'd11060, -25'd8731, 25'd8343, -25'd9605, 25'd8731, 25'd10866, 25'd11254, -25'd10478, 25'd4463}, '{25'd4754, -25'd10381, 25'd3881, -25'd8537, 25'd8634, 25'd485, 25'd7955, -25'd11739, 25'd7276}, '{-25'd6597, 25'd10963, 25'd1649, 25'd7761, -25'd4172, 25'd3105, -25'd2037, 25'd9702, 25'd9411}, '{-25'd5918, 25'd0, -25'd7276, 25'd5821, -25'd4269, -25'd1358, -25'd6403, 25'd1746, 25'd3396}, '{-25'd10090, 25'd11933, -25'd10963, 25'd2425, 25'd6791, 25'd2037, -25'd2134, -25'd3493, 25'd5627}, '{25'd10769, -25'd6403, -25'd10575, 25'd1067, 25'd9799, 25'd8926, -25'd8829, -25'd291, 25'd4075}}, '{'{-25'd8926, 25'd679, 25'd8440, 25'd7082, -25'd7858, -25'd8343, 25'd6403, -25'd9411, 25'd1455}, '{-25'd8829, 25'd11448, 25'd11642, 25'd6791, 25'd10381, 25'd1067, 25'd1843, 25'd12321, -25'd1358}, '{25'd4269, 25'd4075, 25'd7276, -25'd970, -25'd97, -25'd9120, 25'd8731, -25'd4754, -25'd1940}, '{25'd6694, 25'd11642, 25'd10381, -25'd3881, -25'd7470, -25'd10769, 25'd9702, -25'd3396, 25'd11448}, '{-25'd582, 25'd1358, -25'd5045, -25'd970, -25'd4560, -25'd10284, 25'd3590, 25'd10672, -25'd6403}, '{25'd10575, 25'd8537, -25'd2910, -25'd1067, -25'd3008, -25'd6694, -25'd7276, -25'd5918, -25'd6112}, '{25'd4851, -25'd8149, -25'd1455, -25'd11351, 25'd1455, 25'd3105, -25'd1746, -25'd11739, 25'd10187}, '{-25'd1843, 25'd97, -25'd11351, -25'd5627, 25'd582, 25'd5239, -25'd2619, 25'd3396, 25'd1940}, '{25'd2716, -25'd7179, 25'd11642, -25'd9023, 25'd3978, 25'd6403, -25'd11157, -25'd4560, -25'd10769}}, '{'{-25'd8440, 25'd9023, 25'd3105, -25'd8343, -25'd5336, -25'd3299, 25'd7179, 25'd3493, 25'd3493}, '{25'd2328, -25'd970, -25'd8634, -25'd2813, 25'd9411, 25'd12321, -25'd3105, 25'd9605, 25'd6112}, '{25'd7470, 25'd6306, 25'd10381, -25'd8731, 25'd3687, 25'd2813, 25'd4269, -25'd776, 25'd388}, '{-25'd388, -25'd6015, -25'd8829, 25'd11351, 25'd5336, 25'd10478, -25'd6015, -25'd2910, 25'd2231}, '{25'd7470, -25'd9799, -25'd2910, 25'd11448, -25'd4269, -25'd2328, 25'd9702, 25'd7664, 25'd1358}, '{-25'd5336, -25'd7955, -25'd6888, 25'd7082, 25'd12030, 25'd6791, 25'd3978, 25'd1746, 25'd8926}, '{-25'd4269, -25'd7179, -25'd2910, 25'd8634, 25'd6403, -25'd6694, 25'd8343, 25'd873, -25'd5918}, '{-25'd7082, 25'd5142, 25'd5045, -25'd9896, 25'd3396, -25'd7373, 25'd6403, -25'd3202, -25'd2813}, '{-25'd5821, 25'd7567, -25'd5530, 25'd8537, -25'd873, -25'd7761, 25'd6985, -25'd291, -25'd5627}}},
    '{'{'{-25'd204, 25'd6004, 25'd814, -25'd10176, -25'd4477, -25'd9565, -25'd6411, -25'd5088, -25'd1018}, '{25'd8141, -25'd4172, 25'd4274, 25'd12923, -25'd2544, 25'd10990, 25'd4579, 25'd5800, -25'd6309}, '{25'd4172, -25'd9972, -25'd2747, -25'd509, -25'd1832, 25'd10990, 25'd712, 25'd2951, 25'd11193}, '{25'd6716, -25'd611, 25'd305, -25'd6411, -25'd1119, -25'd2747, 25'd10176, -25'd2137, 25'd8548}, '{25'd4681, 25'd1119, -25'd9972, -25'd1526, -25'd9972, 25'd1425, 25'd4884, 25'd7734, 25'd10990}, '{25'd712, -25'd7734, 25'd5393, 25'd10786, -25'd4681, 25'd11092, 25'd1526, 25'd5495, -25'd9463}, '{25'd11804, 25'd7327, 25'd9463, 25'd509, 25'd1425, 25'd6207, -25'd8548, 25'd8751, 25'd6411}, '{-25'd7327, 25'd10176, -25'd7225, 25'd3460, -25'd4376, -25'd1526, -25'd8751, -25'd10176, 25'd3358}, '{25'd6309, 25'd1832, 25'd3765, -25'd5190, 25'd7021, -25'd4681, 25'd712, -25'd6309, -25'd2239}}, '{'{25'd5902, 25'd2646, 25'd7327, -25'd9870, -25'd2646, 25'd3460, 25'd4477, -25'd3867, -25'd9463}, '{-25'd407, 25'd1628, 25'd2442, 25'd8039, 25'd6920, -25'd1119, -25'd12007, -25'd10176, 25'd6614}, '{25'd9667, -25'd712, -25'd3358, 25'd9769, -25'd712, 25'd7225, 25'd3053, 25'd9667, -25'd4172}, '{-25'd8039, 25'd2137, 25'd2646, -25'd6309, -25'd3562, 25'd7937, -25'd4070, 25'd9870, -25'd11804}, '{25'd5698, 25'd8955, -25'd11092, 25'd814, 25'd1221, -25'd2137, -25'd10990, -25'd8141, -25'd5495}, '{-25'd6716, -25'd9565, 25'd2137, 25'd9972, -25'd10481, -25'd3969, 25'd7123, -25'd12821, -25'd9565}, '{25'd2747, -25'd1018, -25'd12007, 25'd9158, 25'd5800, 25'd4884, 25'd7734, -25'd5190, -25'd2137}, '{-25'd9972, 25'd712, -25'd9260, 25'd5902, 25'd7225, 25'd5190, -25'd12414, -25'd4172, -25'd10786}, '{-25'd814, 25'd0, -25'd10074, -25'd407, 25'd5495, 25'd6512, 25'd3358, 25'd2544, -25'd8649}}, '{'{25'd10176, -25'd6818, 25'd9463, -25'd10379, -25'd6614, -25'd9056, 25'd5698, -25'd1221, 25'd9260}, '{25'd4884, -25'd5291, 25'd8242, 25'd916, 25'd3663, 25'd8242, 25'd12618, 25'd509, 25'd6920}, '{25'd7327, -25'd7734, 25'd407, 25'd1425, 25'd2137, 25'd8039, 25'd2951, 25'd7225, -25'd4477}, '{-25'd3562, -25'd611, 25'd7021, 25'd2137, 25'd7734, 25'd6818, 25'd11702, 25'd9972, -25'd5800}, '{25'd5800, 25'd10583, 25'd7327, -25'd204, -25'd2544, 25'd4376, -25'd814, -25'd7225, -25'd9463}, '{25'd6716, -25'd916, 25'd4884, 25'd9565, 25'd8446, -25'd10481, -25'd3256, 25'd6512, 25'd10481}, '{25'd10583, 25'd7632, 25'd2544, 25'd814, -25'd2340, 25'd2747, -25'd2747, 25'd10786, 25'd5800}, '{-25'd1323, 25'd9972, 25'd2951, -25'd7632, -25'd6512, -25'd5291, 25'd7123, 25'd6309, 25'd7835}, '{25'd4681, -25'd2442, -25'd7327, 25'd9870, 25'd4783, 25'd6512, 25'd8344, 25'd3969, -25'd4376}}},
    '{'{'{25'd425, -25'd6804, 25'd7123, -25'd4146, -25'd1595, -25'd2870, 25'd11163, 25'd7017, 25'd11057}, '{25'd4253, 25'd3508, -25'd8930, -25'd5847, -25'd9674, 25'd5635, 25'd2764, 25'd851, 25'd957}, '{25'd12013, 25'd638, 25'd7655, -25'd9781, 25'd9462, 25'd9037, -25'd7655, 25'd3615, 25'd5209}, '{25'd13289, 25'd5954, 25'd9781, -25'd9143, 25'd2126, -25'd3083, 25'd8824, 25'd7761, 25'd11269}, '{-25'd1063, -25'd8292, 25'd12864, -25'd4678, 25'd3721, -25'd6485, -25'd1914, 25'd5103, -25'd2339}, '{-25'd3721, 25'd11057, 25'd4359, 25'd8930, 25'd2658, -25'd7123, 25'd1063, 25'd425, -25'd7655}, '{25'd11375, -25'd5209, 25'd8292, -25'd1488, -25'd4678, -25'd4678, 25'd4359, -25'd5316, -25'd10100}, '{-25'd5847, 25'd4359, 25'd3615, -25'd8080, 25'd1595, -25'd5103, 25'd9674, -25'd4890, -25'd851}, '{-25'd8505, -25'd7229, 25'd12120, 25'd10950, 25'd11269, 25'd2445, 25'd1701, -25'd9037, -25'd2764}}, '{'{-25'd8080, -25'd4890, -25'd9356, 25'd6910, -25'd12013, -25'd5209, 25'd2126, 25'd7123, -25'd5741}, '{-25'd4678, -25'd2233, 25'd5741, -25'd1701, 25'd9143, -25'd3083, -25'd8505, 25'd4040, -25'd4571}, '{25'd3296, -25'd12013, 25'd0, 25'd3296, -25'd6698, -25'd9887, 25'd4253, -25'd3189, -25'd5316}, '{-25'd2764, -25'd5316, 25'd10100, -25'd10206, -25'd11163, -25'd8505, -25'd3827, -25'd5316, -25'd6379}, '{25'd8399, -25'd13502, 25'd6698, -25'd2020, -25'd3083, 25'd5209, -25'd5847, -25'd4146, 25'd744}, '{-25'd9887, -25'd6804, 25'd6910, 25'd9462, -25'd10419, -25'd4253, 25'd8505, -25'd638, 25'd3083}, '{25'd5422, 25'd7761, 25'd1595, -25'd12013, -25'd7867, 25'd7336, 25'd9249, -25'd10950, 25'd5847}, '{-25'd5954, -25'd1063, -25'd3189, -25'd10950, -25'd5316, 25'd2126, 25'd3083, -25'd12651, 25'd2870}, '{-25'd9568, -25'd9781, 25'd6166, -25'd2764, 25'd6485, -25'd8611, 25'd9993, 25'd1488, 25'd2764}}, '{'{25'd3083, -25'd9674, 25'd7761, 25'd8186, -25'd3827, -25'd5635, 25'd10738, 25'd13289, 25'd13076}, '{25'd10738, -25'd3508, 25'd1276, 25'd6060, 25'd9356, 25'd8505, -25'd5209, -25'd5316, 25'd213}, '{25'd7017, 25'd9674, -25'd1488, -25'd9993, -25'd2977, 25'd13289, 25'd3827, 25'd12226, -25'd4784}, '{25'd11588, -25'd1488, -25'd6804, 25'd2764, 25'd12439, 25'd6379, -25'd6272, -25'd6804, -25'd3402}, '{25'd11694, 25'd2764, -25'd9356, 25'd9674, -25'd6910, 25'd10206, -25'd5741, -25'd7229, -25'd2233}, '{-25'd10100, 25'd0, -25'd957, 25'd6379, 25'd11801, 25'd9993, -25'd6591, 25'd425, 25'd9993}, '{25'd11588, -25'd9568, 25'd7655, 25'd11694, 25'd8186, 25'd744, -25'd4146, 25'd2126, -25'd4678}, '{25'd1488, 25'd1595, 25'd6485, 25'd8718, 25'd8399, 25'd6272, 25'd10419, -25'd4571, 25'd4253}, '{25'd319, 25'd7867, -25'd1807, 25'd9568, 25'd7867, -25'd3402, -25'd6166, -25'd2764, -25'd3827}}},
    '{'{'{25'd1127, 25'd7516, 25'd0, 25'd6890, 25'd501, -25'd877, -25'd752, 25'd0, 25'd4760}, '{-25'd3132, 25'd125, 25'd7015, 25'd5261, -25'd1378, -25'd3633, -25'd4635, 25'd2505, -25'd8518}, '{-25'd5011, 25'd6890, -25'd1002, 25'd10272, 25'd1127, 25'd4510, -25'd10146, -25'd5762, -25'd1879}, '{-25'd6639, 25'd9896, 25'd376, -25'd1127, -25'd9019, -25'd10021, 25'd8518, 25'd11775, -25'd1628}, '{-25'd10021, -25'd9645, -25'd7641, -25'd3883, 25'd12526, 25'd12151, -25'd9896, 25'd12151, 25'd10146}, '{25'd8267, 25'd10146, 25'd11149, -25'd1253, 25'd10146, -25'd9520, 25'd11399, -25'd2505, -25'd3758}, '{-25'd5386, 25'd10522, 25'd1879, -25'd2129, 25'd10522, 25'd14531, 25'd11775, 25'd2631, 25'd125}, '{-25'd7391, -25'd4134, -25'd1503, -25'd6388, 25'd10522, 25'd8643, 25'd1879, 25'd2004, 25'd1754}, '{-25'd8267, 25'd7516, 25'd11900, -25'd5762, 25'd2631, -25'd4259, -25'd4134, 25'd4510, 25'd13403}}, '{'{25'd15909, 25'd4760, -25'd6013, -25'd5261, 25'd8768, -25'd4760, 25'd2756, -25'd5386, -25'd3382}, '{25'd376, 25'd7516, 25'd9645, -25'd2881, -25'd2129, 25'd8518, 25'd6764, -25'd7641, -25'd12151}, '{-25'd5887, -25'd12276, 25'd5762, 25'd7516, -25'd1628, -25'd1002, -25'd10146, 25'd4008, -25'd8393}, '{25'd11023, -25'd9144, 25'd3006, -25'd10773, 25'd8267, 25'd5136, 25'd6514, 25'd9270, -25'd11023}, '{25'd5136, -25'd2505, -25'd5261, 25'd9019, -25'd501, 25'd9019, -25'd8393, 25'd3132, -25'd1879}, '{25'd7516, -25'd3006, -25'd3507, -25'd7766, 25'd5136, 25'd5386, -25'd2505, -25'd11524, 25'd1628}, '{-25'd12276, -25'd877, -25'd7641, 25'd2756, -25'd12526, -25'd4008, -25'd3633, -25'd1002, -25'd9645}, '{25'd5386, -25'd10773, 25'd5386, -25'd8017, -25'd6013, 25'd4760, 25'd9520, -25'd7641, 25'd1127}, '{-25'd6890, -25'd14030, 25'd7641, -25'd5011, -25'd6388, 25'd3257, -25'd125, -25'd5261, 25'd5512}}, '{'{25'd877, -25'd6639, -25'd6013, -25'd2255, -25'd4635, -25'd2255, -25'd4885, 25'd6138, -25'd4635}, '{25'd501, 25'd9395, -25'd4134, 25'd9019, -25'd2004, 25'd12151, 25'd5762, -25'd4760, 25'd4134}, '{25'd9520, 25'd6263, 25'd10522, 25'd12276, 25'd10021, -25'd6764, -25'd376, -25'd1628, -25'd7140}, '{-25'd4510, 25'd3006, -25'd1754, -25'd2255, -25'd752, 25'd11399, -25'd6263, -25'd3382, -25'd8518}, '{-25'd2505, 25'd4885, 25'd2255, 25'd9395, -25'd6890, 25'd6764, -25'd5512, -25'd2255, 25'd10146}, '{25'd11524, -25'd9645, -25'd9019, -25'd1253, -25'd3257, -25'd7892, 25'd1127, -25'd4510, -25'd6514}, '{-25'd4384, 25'd3006, 25'd626, 25'd1253, -25'd6013, -25'd5762, 25'd3257, 25'd5386, -25'd3257}, '{-25'd11399, 25'd4134, 25'd3883, -25'd10272, 25'd7391, 25'd4384, -25'd251, 25'd1378, -25'd8142}, '{25'd2505, -25'd2004, 25'd4259, -25'd4760, 25'd10397, 25'd4384, -25'd6639, 25'd9771, -25'd7265}}},
    '{'{'{25'd2827, -25'd7324, -25'd11821, 25'd128, -25'd4112, -25'd2313, -25'd12463, -25'd13748, -25'd3726}, '{25'd2441, -25'd3469, 25'd4497, -25'd10022, 25'd5782, -25'd2570, 25'd2056, -25'd13491, -25'd8480}, '{-25'd5397, -25'd5140, 25'd8609, 25'd4369, -25'd3341, 25'd2570, 25'd2184, 25'd385, -25'd12078}, '{25'd6039, -25'd4754, 25'd7709, 25'd1927, -25'd2441, -25'd10793, -25'd1285, -25'd2056, -25'd7581}, '{-25'd7966, 25'd1285, 25'd2955, 25'd3983, 25'd5140, -25'd8095, -25'd2056, 25'd5910, -25'd8609}, '{-25'd3983, 25'd2698, 25'd11179, 25'd8866, 25'd3598, -25'd10665, -25'd2441, -25'd8866, 25'd10022}, '{-25'd7195, -25'd11050, 25'd11435, 25'd2570, 25'd12335, 25'd257, -25'd3726, -25'd9380, 25'd4754}, '{-25'd7581, -25'd642, 25'd5140, 25'd6424, 25'd9123, 25'd2698, -25'd3212, 25'd8480, -25'd9251}, '{25'd7067, 25'd7324, 25'd9765, -25'd1285, 25'd3598, 25'd2570, -25'd10793, 25'd9508, 25'd1413}}, '{'{-25'd9251, -25'd6039, -25'd2570, 25'd9251, 25'd899, 25'd4112, -25'd10922, 25'd2570, -25'd10408}, '{-25'd2441, -25'd4626, 25'd7581, 25'd10536, 25'd8994, 25'd3469, -25'd16447, -25'd6553, -25'd6167}, '{25'd11050, -25'd2698, 25'd6938, -25'd11949, -25'd2441, 25'd3469, 25'd7195, -25'd1028, -25'd2441}, '{-25'd8095, -25'd6810, 25'd6938, -25'd10151, 25'd1927, -25'd11692, 25'd3341, 25'd3341, 25'd4369}, '{25'd2184, -25'd9637, 25'd4369, 25'd4112, 25'd7966, -25'd1799, 25'd2056, -25'd4754, -25'd2184}, '{25'd3855, 25'd1927, -25'd257, -25'd9508, -25'd11179, -25'd1799, -25'd4883, 25'd7966, -25'd10536}, '{25'd1285, -25'd128, -25'd12206, 25'd771, 25'd5654, -25'd1285, 25'd5782, 25'd1285, 25'd2184}, '{-25'd1799, -25'd13748, 25'd2827, 25'd4240, -25'd10151, -25'd514, -25'd11692, -25'd3469, 25'd771}, '{-25'd3598, 25'd5397, 25'd1413, 25'd9251, 25'd8095, -25'd12335, 25'd2698, -25'd7581, 25'd7581}}, '{'{-25'd9508, -25'd9765, -25'd2570, -25'd8480, 25'd3341, 25'd7195, -25'd3855, -25'd10536, 25'd1156}, '{-25'd1028, -25'd12592, 25'd13877, -25'd2955, 25'd7838, -25'd4240, -25'd9508, -25'd7195, -25'd10151}, '{25'd771, 25'd7966, 25'd10922, 25'd4112, 25'd6938, 25'd7709, 25'd8352, 25'd2313, -25'd642}, '{-25'd2827, 25'd9765, 25'd15290, 25'd385, 25'd14648, 25'd1156, 25'd4240, -25'd10536, -25'd3855}, '{25'd9765, -25'd8609, -25'd3084, 25'd7195, 25'd2955, -25'd6296, 25'd8609, -25'd4112, 25'd2056}, '{-25'd1285, -25'd1799, -25'd771, 25'd5140, -25'd128, -25'd4497, 25'd5140, 25'd5268, 25'd9380}, '{-25'd385, 25'd8866, 25'd2184, 25'd3726, 25'd11692, 25'd12078, 25'd11050, 25'd4240, 25'd7709}, '{25'd7452, 25'd14262, -25'd2827, -25'd2056, -25'd6553, 25'd5140, 25'd10536, 25'd2056, -25'd6296}, '{25'd12078, -25'd1927, 25'd7838, -25'd5011, 25'd13363, 25'd14005, 25'd5782, 25'd6681, -25'd3084}}},
    '{'{'{25'd3489, -25'd9091, -25'd2326, -25'd9408, -25'd3700, -25'd9620, 25'd8246, -25'd11734, 25'd3066}, '{25'd9620, 25'd10888, 25'd1480, 25'd951, 25'd8563, 25'd10677, 25'd3171, 25'd11840, -25'd7717}, '{-25'd8668, 25'd5920, 25'd3066, -25'd5391, -25'd5180, 25'd9514, 25'd9303, 25'd11945, 25'd7506}, '{-25'd7823, 25'd6871, -25'd5180, 25'd423, 25'd9620, -25'd6131, 25'd3806, 25'd529, -25'd2854}, '{25'd7717, -25'd2537, -25'd9937, 25'd106, -25'd5391, -25'd2114, 25'd12474, -25'd8563, -25'd1480}, '{25'd7823, 25'd7928, -25'd10360, -25'd8668, 25'd634, 25'd5814, -25'd8351, 25'd5074, 25'd8563}, '{-25'd3383, -25'd10888, 25'd10571, 25'd2960, 25'd6343, 25'd7083, 25'd7188, 25'd106, 25'd8034}, '{25'd4863, 25'd11206, -25'd7611, -25'd5603, -25'd211, 25'd9408, -25'd2854, 25'd6660, 25'd7188}, '{-25'd5814, 25'd4968, 25'd7506, -25'd6343, 25'd6237, 25'd7188, 25'd8351, 25'd5603, -25'd10783}}, '{'{-25'd423, -25'd846, -25'd13531, -25'd6977, -25'd5603, -25'd12580, 25'd1586, 25'd3594, 25'd4228}, '{-25'd740, 25'd5286, 25'd5708, -25'd9091, -25'd8351, 25'd9726, -25'd4123, 25'd1269, -25'd4651}, '{25'd6554, 25'd9831, 25'd10043, -25'd5286, -25'd5920, -25'd3806, -25'd2431, 25'd6660, 25'd8246}, '{-25'd2854, -25'd10466, -25'd10254, 25'd9831, -25'd1480, 25'd4863, -25'd2220, 25'd7928, 25'd3911}, '{25'd8774, 25'd3806, -25'd7188, -25'd3383, -25'd6237, 25'd9408, 25'd2854, 25'd12791, -25'd4334}, '{-25'd634, 25'd5391, -25'd7294, -25'd10043, -25'd8668, -25'd9303, -25'd1163, -25'd7928, -25'd2537}, '{-25'd1903, 25'd5603, 25'd6026, -25'd11523, 25'd4440, 25'd3911, 25'd423, 25'd5603, 25'd8668}, '{-25'd9726, 25'd8880, 25'd10148, -25'd2220, -25'd3277, -25'd529, 25'd8140, 25'd2114, -25'd529}, '{25'd3700, -25'd7717, 25'd8140, -25'd634, 25'd2220, 25'd3383, -25'd4440, 25'd5708, -25'd7823}}, '{'{-25'd12897, -25'd5074, 25'd7928, -25'd12791, -25'd11840, 25'd6026, -25'd9620, -25'd8563, 25'd2749}, '{25'd4228, -25'd11840, -25'd6871, 25'd10571, 25'd4546, 25'd5708, 25'd8140, 25'd9726, 25'd8140}, '{-25'd10466, -25'd10994, 25'd3277, 25'd5286, -25'd8880, 25'd5920, 25'd11100, -25'd9197, 25'd5920}, '{25'd5286, 25'd11945, 25'd634, 25'd529, -25'd8880, 25'd8457, 25'd8246, 25'd3383, 25'd4228}, '{25'd9197, -25'd4017, 25'd10466, 25'd1057, -25'd4334, -25'd7294, 25'd12368, -25'd8246, -25'd8668}, '{25'd8668, -25'd9620, -25'd10571, 25'd3806, 25'd0, 25'd7928, -25'd7294, 25'd8986, 25'd423}, '{-25'd10783, 25'd1903, -25'd106, -25'd951, -25'd10677, -25'd3911, 25'd529, -25'd3171, -25'd7611}, '{25'd7506, -25'd9091, -25'd3700, 25'd3277, 25'd6237, 25'd2643, 25'd10783, -25'd1480, -25'd3383}, '{-25'd3911, -25'd8034, -25'd10783, 25'd11206, 25'd3806, 25'd9726, 25'd7611, -25'd10360, -25'd2114}}},
    '{'{'{-25'd11634, -25'd7168, 25'd470, 25'd6228, 25'd5406, -25'd13867, 25'd7638, -25'd5288, 25'd13632}, '{-25'd12457, -25'd1293, -25'd353, -25'd11164, 25'd4818, -25'd470, -25'd11986, 25'd9636, 25'd9401}, '{25'd1293, -25'd4231, 25'd8108, -25'd10106, -25'd11634, 25'd6698, 25'd3643, 25'd235, 25'd235}, '{25'd6581, -25'd11751, -25'd4583, 25'd2350, -25'd10224, -25'd12927, -25'd4231, 25'd1880, 25'd12692}, '{-25'd11516, 25'd6228, -25'd3525, -25'd5053, -25'd13867, -25'd5523, -25'd7168, 25'd4348, 25'd12809}, '{-25'd1058, 25'd3525, 25'd2350, 25'd3995, 25'd8344, 25'd2703, -25'd12574, 25'd12104, -25'd470}, '{-25'd353, 25'd5406, -25'd13984, -25'd3408, 25'd1175, 25'd8814, 25'd8579, -25'd6933, 25'd11516}, '{-25'd11281, -25'd470, 25'd5641, 25'd3525, -25'd2115, 25'd2703, 25'd4583, -25'd5523, 25'd13632}, '{25'd2938, 25'd7403, 25'd4701, -25'd5758, -25'd7521, -25'd3408, -25'd1058, 25'd14924, 25'd7756}}, '{'{-25'd8461, 25'd3643, 25'd7168, 25'd118, -25'd6933, -25'd7756, -25'd7991, -25'd5993, 25'd9401}, '{-25'd9871, -25'd7873, 25'd12104, -25'd8579, 25'd2820, 25'd3173, -25'd9519, 25'd1293, 25'd5523}, '{25'd9636, 25'd10106, 25'd1763, 25'd8344, 25'd10459, -25'd11634, 25'd6111, 25'd3290, -25'd5641}, '{-25'd235, -25'd9049, 25'd3408, 25'd2468, -25'd5993, 25'd7403, -25'd9166, -25'd5171, -25'd2820}, '{25'd7521, 25'd7403, -25'd8461, -25'd10929, -25'd5406, 25'd353, 25'd235, 25'd118, -25'd4701}, '{-25'd8461, -25'd3760, 25'd3878, -25'd353, 25'd2233, -25'd13044, -25'd1293, -25'd7521, 25'd4231}, '{-25'd7756, -25'd11869, -25'd940, 25'd2350, -25'd2820, 25'd5993, -25'd7638, 25'd0, 25'd235}, '{25'd5876, -25'd7638, 25'd1293, -25'd11986, -25'd10929, 25'd9519, -25'd470, 25'd9166, 25'd7756}, '{25'd4348, 25'd9989, 25'd5641, 25'd6933, 25'd11281, 25'd2468, -25'd4113, 25'd12809, 25'd12222}}, '{'{-25'd7991, 25'd6698, 25'd5641, -25'd7873, -25'd6816, -25'd8696, -25'd2938, -25'd940, -25'd11869}, '{25'd9049, -25'd2350, -25'd940, -25'd1058, 25'd3995, 25'd7638, 25'd1058, 25'd10224, -25'd11869}, '{-25'd7873, 25'd8931, 25'd1998, -25'd7286, 25'd1880, 25'd1058, -25'd6228, 25'd3878, 25'd1645}, '{-25'd9284, 25'd2115, 25'd9636, -25'd6463, -25'd4113, 25'd5053, 25'd1175, 25'd3995, 25'd2115}, '{-25'd1410, -25'd6698, -25'd11281, 25'd1645, -25'd7168, 25'd9519, -25'd8579, -25'd2820, 25'd7756}, '{25'd2938, -25'd8344, -25'd3173, 25'd5876, 25'd5053, -25'd1528, -25'd10341, -25'd9166, -25'd9636}, '{25'd8108, -25'd12457, 25'd6698, 25'd7286, -25'd4113, -25'd8226, -25'd7756, 25'd588, 25'd10811}, '{-25'd5171, 25'd4818, -25'd2703, -25'd5523, -25'd10811, -25'd10224, -25'd1175, 25'd6463, 25'd13514}, '{25'd470, -25'd5758, 25'd1998, 25'd588, 25'd8108, -25'd5171, -25'd4936, -25'd9284, -25'd2820}}},
    '{'{'{25'd8739, -25'd3440, -25'd7438, 25'd2789, -25'd7438, 25'd3719, 25'd1859, -25'd6973, -25'd2138}, '{25'd8274, 25'd5857, -25'd1952, -25'd2138, 25'd9018, -25'd2417, -25'd8089, 25'd5950, -25'd5950}, '{-25'd5578, -25'd3998, -25'd8739, -25'd2789, 25'd10692, 25'd186, -25'd5485, -25'd5020, -25'd6322}, '{25'd744, 25'd3347, 25'd10227, 25'd4742, 25'd1209, 25'd9018, -25'd5950, 25'd4277, 25'd7624}, '{-25'd7159, -25'd3719, 25'd9948, 25'd9111, -25'd9204, -25'd5299, 25'd2138, -25'd1766, 25'd10041}, '{25'd5299, -25'd6322, 25'd9762, 25'd1023, -25'd3905, -25'd7438, 25'd372, -25'd4370, -25'd6508}, '{25'd4463, 25'd186, -25'd3161, -25'd10134, 25'd837, 25'd2510, 25'd0, 25'd8739, 25'd6043}, '{25'd5485, 25'd9204, 25'd10506, 25'd1023, -25'd10506, 25'd6508, -25'd1488, -25'd1302, -25'd1859}, '{-25'd9390, -25'd1581, 25'd651, -25'd3998, 25'd6415, 25'd9762, 25'd10878, 25'd6973, -25'd6694}}, '{'{-25'd2975, 25'd8739, -25'd5299, -25'd7996, 25'd9576, -25'd2417, 25'd1116, 25'd6322, 25'd1302}, '{25'd3533, -25'd372, 25'd4835, 25'd5485, -25'd3626, -25'd1209, -25'd2417, 25'd7810, 25'd5299}, '{25'd465, -25'd3068, -25'd11157, -25'd93, 25'd9297, 25'd1859, -25'd7810, -25'd2324, 25'd10878}, '{25'd11435, -25'd7345, -25'd5020, 25'd7252, -25'd4742, 25'd7996, -25'd9855, 25'd9204, -25'd5299}, '{25'd5392, 25'd3068, -25'd7531, 25'd3254, 25'd11064, 25'd5671, -25'd3812, 25'd8646, -25'd4091}, '{-25'd9111, -25'd7531, 25'd1302, -25'd5764, -25'd2231, -25'd7531, 25'd6136, 25'd5950, 25'd3812}, '{25'd8089, 25'd9390, -25'd8181, 25'd186, 25'd4835, -25'd5671, -25'd3347, -25'd10041, -25'd1395}, '{25'd8367, -25'd3347, 25'd4277, -25'd5578, 25'd3440, 25'd11250, -25'd2882, -25'd6880, -25'd8832}, '{25'd10971, 25'd7066, -25'd6043, -25'd9576, 25'd8739, 25'd8460, -25'd8646, 25'd5020, -25'd6322}}, '{'{-25'd7810, 25'd651, 25'd1116, -25'd4463, 25'd3812, 25'd9018, 25'd1116, 25'd5206, -25'd2789}, '{-25'd8739, 25'd2510, 25'd10506, 25'd10971, 25'd1673, 25'd1116, 25'd3998, 25'd6043, 25'd2231}, '{-25'd10785, -25'd9018, -25'd7345, 25'd10971, -25'd9018, -25'd279, 25'd3068, -25'd11900, 25'd11064}, '{-25'd10041, 25'd9390, -25'd2510, -25'd10506, -25'd1581, -25'd2789, -25'd558, 25'd1302, -25'd5206}, '{25'd2789, 25'd5299, 25'd744, 25'd5764, 25'd372, -25'd7252, 25'd3812, 25'd2045, -25'd3533}, '{-25'd1673, 25'd3347, -25'd6229, -25'd10599, 25'd9948, -25'd651, 25'd7159, 25'd7717, 25'd6601}, '{-25'd10227, 25'd2510, 25'd3905, 25'd3068, 25'd558, 25'd2324, 25'd0, 25'd10134, -25'd9576}, '{-25'd4835, 25'd186, -25'd9483, -25'd7624, 25'd8089, -25'd8460, 25'd4927, 25'd6136, 25'd2789}, '{25'd3347, 25'd465, 25'd2510, -25'd1673, -25'd1023, -25'd9204, -25'd2138, 25'd8553, -25'd6229}}},
    '{'{'{-25'd9728, 25'd9011, 25'd0, 25'd4915, 25'd6451, 25'd512, 25'd3277, 25'd6349, 25'd7066}, '{-25'd614, 25'd307, -25'd2662, -25'd9216, 25'd5530, 25'd3686, -25'd3584, 25'd7578, 25'd6656}, '{-25'd4198, -25'd10854, 25'd5222, -25'd1024, 25'd5530, -25'd6758, 25'd10752, -25'd4096, -25'd2355}, '{25'd11366, -25'd6758, -25'd2867, -25'd205, -25'd9421, -25'd5632, 25'd410, -25'd12083, 25'd3072}, '{-25'd5120, 25'd4710, 25'd5325, 25'd1843, 25'd9626, -25'd1843, -25'd3174, -25'd2355, 25'd2150}, '{25'd3277, -25'd8602, -25'd1331, 25'd5018, 25'd2867, -25'd5222, -25'd13005, 25'd5018, -25'd10957}, '{-25'd6656, 25'd8602, 25'd1126, 25'd3994, -25'd3686, -25'd6963, 25'd7782, 25'd8192, -25'd6963}, '{25'd6554, -25'd5325, 25'd7680, 25'd8090, 25'd8294, -25'd10035, -25'd11264, 25'd3482, -25'd1536}, '{25'd7578, -25'd1229, 25'd7680, 25'd3379, 25'd6246, -25'd7680, -25'd11366, -25'd1536, -25'd410}}, '{'{25'd9830, 25'd7475, 25'd11776, -25'd5837, 25'd4813, 25'd13005, -25'd3072, -25'd717, 25'd614}, '{-25'd3891, 25'd1741, 25'd12902, 25'd3482, 25'd4506, 25'd11776, -25'd6144, 25'd922, -25'd1946}, '{25'd6042, -25'd2048, 25'd9626, -25'd819, -25'd9523, -25'd9216, -25'd5734, 25'd5120, -25'd1536}, '{25'd11469, -25'd7578, -25'd4915, 25'd7475, 25'd3584, -25'd4915, -25'd1024, -25'd4403, -25'd3891}, '{25'd4403, -25'd410, -25'd1741, 25'd3379, -25'd10854, 25'd9216, -25'd1843, -25'd1946, -25'd9523}, '{-25'd8294, 25'd3379, -25'd3379, 25'd11162, 25'd7066, -25'd6656, 25'd2355, -25'd10854, 25'd8499}, '{25'd11981, 25'd2560, 25'd717, -25'd5837, 25'd5222, 25'd1434, -25'd2150, -25'd5734, 25'd102}, '{25'd2355, 25'd2560, 25'd11469, 25'd9318, 25'd3277, -25'd102, -25'd307, 25'd10035, 25'd7885}, '{-25'd8397, 25'd614, -25'd410, -25'd5427, 25'd2253, 25'd6451, 25'd4096, 25'd2560, -25'd4710}}, '{'{25'd2867, -25'd614, 25'd5939, 25'd8602, -25'd10650, -25'd10240, 25'd2662, 25'd102, -25'd7680}, '{25'd1229, -25'd1946, -25'd3072, 25'd205, -25'd6451, -25'd2560, 25'd4608, -25'd7885, 25'd5837}, '{25'd9318, -25'd9318, 25'd1126, 25'd9830, -25'd3174, 25'd5018, -25'd10854, 25'd9421, 25'd8499}, '{25'd4813, -25'd8806, 25'd1331, 25'd205, 25'd8909, 25'd1229, -25'd2253, 25'd1638, 25'd2867}, '{-25'd1946, -25'd4096, -25'd8806, -25'd1126, -25'd3482, -25'd3379, 25'd4198, -25'd12083, 25'd8602}, '{-25'd6144, -25'd410, -25'd1024, -25'd2150, -25'd4301, 25'd6349, 25'd2355, -25'd11366, 25'd6144}, '{25'd8192, -25'd2662, 25'd12186, 25'd7782, -25'd819, -25'd5632, 25'd2253, -25'd10445, 25'd5939}, '{-25'd1638, -25'd5120, -25'd4915, 25'd1024, 25'd922, 25'd1331, -25'd4813, -25'd2662, 25'd9421}, '{25'd1536, -25'd6451, 25'd2662, 25'd10240, -25'd6349, 25'd7066, 25'd7987, -25'd6451, 25'd2150}}},
    '{'{'{25'd3960, 25'd8602, 25'd5052, 25'd2867, 25'd11743, 25'd8602, -25'd7374, 25'd2321, -25'd5325}, '{-25'd7920, -25'd9558, -25'd4506, -25'd9012, 25'd10924, -25'd1775, 25'd9968, -25'd8739, -25'd3823}, '{25'd12153, -25'd4096, 25'd10787, 25'd5325, 25'd3960, 25'd12016, 25'd6418, 25'd2048, 25'd7920}, '{25'd5598, -25'd9558, -25'd7374, 25'd5872, 25'd14064, 25'd410, -25'd2048, 25'd8739, 25'd13245}, '{25'd6008, 25'd13655, 25'd13382, 25'd13928, 25'd7100, -25'd6691, -25'd1502, 25'd15430, 25'd546}, '{-25'd6008, -25'd3414, 25'd4096, -25'd273, 25'd3141, -25'd8193, 25'd273, 25'd3414, 25'd8466}, '{-25'd1365, 25'd12289, 25'd9558, 25'd13791, 25'd8739, 25'd13928, 25'd15430, -25'd3004, 25'd11880}, '{-25'd10924, 25'd9149, -25'd2731, 25'd14201, 25'd13655, 25'd6008, 25'd11197, -25'd3550, 25'd14064}, '{25'd1502, 25'd1912, -25'd6691, 25'd8193, 25'd1365, -25'd5735, 25'd11470, -25'd6554, -25'd4233}}, '{'{25'd3414, -25'd2458, -25'd3687, -25'd5872, -25'd12016, -25'd1365, 25'd956, 25'd683, -25'd410}, '{-25'd3141, -25'd12562, 25'd7783, -25'd10651, -25'd12562, 25'd6827, -25'd9285, -25'd1229, -25'd1229}, '{25'd6554, -25'd1365, -25'd7647, -25'd819, -25'd15157, -25'd7100, -25'd15976, 25'd2185, -25'd16249}, '{-25'd12289, -25'd1639, -25'd10378, -25'd5462, -25'd2594, -25'd8056, -25'd14884, -25'd14747, 25'd6418}, '{25'd6964, -25'd10651, 25'd4779, -25'd16659, -25'd9831, -25'd2321, -25'd6008, -25'd4096, -25'd10241}, '{-25'd15430, -25'd7510, -25'd4779, 25'd2048, -25'd9422, -25'd410, -25'd16386, -25'd5052, -25'd9012}, '{25'd819, 25'd5052, -25'd16249, -25'd8739, 25'd2185, -25'd15566, -25'd12426, -25'd14337, -25'd956}, '{25'd1775, -25'd9968, -25'd13245, -25'd17341, 25'd4506, -25'd14884, -25'd12835, -25'd10924, -25'd15703}, '{25'd3004, 25'd3004, -25'd2321, 25'd2048, -25'd6964, -25'd2321, -25'd10104, -25'd14064, 25'd1639}}, '{'{-25'd9149, 25'd683, 25'd5189, 25'd2321, -25'd3414, -25'd1912, -25'd956, 25'd12562, 25'd3414}, '{-25'd2048, 25'd5872, 25'd10924, 25'd11606, 25'd8466, 25'd6691, 25'd8466, 25'd13655, -25'd5872}, '{-25'd1365, -25'd9149, 25'd6008, -25'd5872, 25'd6827, -25'd5052, 25'd5325, 25'd13245, -25'd683}, '{25'd4779, 25'd11606, -25'd4779, -25'd6964, 25'd7100, 25'd3550, -25'd1912, 25'd7510, 25'd10514}, '{25'd3141, -25'd2594, -25'd4096, -25'd6008, 25'd8193, -25'd7920, 25'd9422, -25'd7100, -25'd7783}, '{25'd6281, 25'd9012, 25'd11470, 25'd5325, -25'd1092, -25'd6008, 25'd9695, -25'd5735, 25'd4506}, '{25'd11606, 25'd3960, -25'd7374, -25'd7783, 25'd819, 25'd8056, -25'd4643, 25'd7100, 25'd11333}, '{25'd7100, 25'd0, -25'd9012, -25'd2048, -25'd3687, -25'd8602, 25'd137, -25'd4096, 25'd4369}, '{-25'd4506, 25'd4369, 25'd10514, -25'd8602, -25'd3550, 25'd5462, -25'd4779, 25'd10241, -25'd9012}}},
    '{'{'{25'd7737, -25'd4999, -25'd3809, -25'd12022, -25'd2738, 25'd5118, -25'd1071, 25'd6071, 25'd5714}, '{-25'd119, -25'd12141, -25'd5237, -25'd12499, -25'd13332, -25'd4523, 25'd8213, -25'd2738, 25'd2976}, '{-25'd11427, 25'd5476, 25'd4285, -25'd10832, -25'd15117, -25'd6428, 25'd2500, 25'd3690, 25'd4761}, '{-25'd4999, 25'd4523, -25'd4404, 25'd5476, 25'd6309, -25'd13689, 25'd2857, -25'd10237, -25'd9285}, '{-25'd2500, -25'd3095, -25'd1309, -25'd4285, -25'd3928, -25'd7261, 25'd10356, 25'd10832, -25'd2381}, '{-25'd9285, -25'd7499, -25'd7261, -25'd119, -25'd11308, 25'd1905, -25'd1666, 25'd10594, 25'd9880}, '{25'd119, 25'd9047, -25'd6309, -25'd2262, -25'd7142, 25'd8213, -25'd1071, -25'd8213, 25'd5952}, '{-25'd714, -25'd1547, -25'd714, 25'd7975, -25'd2262, 25'd7618, 25'd5118, 25'd11308, 25'd14046}, '{25'd2619, 25'd10356, 25'd5595, 25'd5118, 25'd9404, 25'd12022, 25'd3809, 25'd2024, -25'd6666}}, '{'{25'd952, -25'd6547, 25'd0, 25'd8094, 25'd9642, 25'd6428, -25'd7380, 25'd1786, 25'd5833}, '{25'd4047, 25'd2738, -25'd1547, -25'd9999, 25'd238, -25'd12856, 25'd8213, 25'd10237, 25'd8809}, '{25'd3095, 25'd1190, -25'd13094, -25'd357, -25'd6904, 25'd6547, -25'd10118, -25'd3928, -25'd9404}, '{25'd6428, -25'd7737, 25'd6071, -25'd9404, -25'd13094, 25'd2500, 25'd11784, -25'd4642, 25'd2024}, '{25'd12022, -25'd6666, -25'd11665, -25'd2738, 25'd11546, 25'd10475, 25'd8928, 25'd4642, -25'd2143}, '{25'd8809, -25'd1428, 25'd7618, 25'd1666, -25'd9523, -25'd9166, 25'd8570, -25'd1786, 25'd9166}, '{-25'd3928, 25'd0, -25'd10118, 25'd10475, -25'd3690, 25'd9999, 25'd1309, -25'd7380, -25'd5595}, '{25'd7737, -25'd3571, 25'd4047, 25'd6547, 25'd6428, 25'd1309, -25'd952, -25'd1666, -25'd1547}, '{-25'd8809, 25'd1666, -25'd3095, -25'd8451, 25'd8809, -25'd10713, -25'd1428, 25'd10356, -25'd8570}}, '{'{25'd11427, 25'd5595, -25'd357, -25'd11665, 25'd4642, 25'd12022, -25'd1190, 25'd357, 25'd12022}, '{25'd357, -25'd1428, 25'd10475, -25'd6190, -25'd1547, 25'd6071, -25'd1666, -25'd7142, 25'd1666}, '{25'd1309, -25'd11070, -25'd12260, -25'd11546, 25'd5118, 25'd11784, -25'd5595, -25'd7856, -25'd2262}, '{25'd7618, 25'd8213, 25'd8094, -25'd6428, 25'd8332, 25'd357, -25'd9880, 25'd11784, -25'd5237}, '{25'd2143, -25'd2143, 25'd11189, 25'd8094, -25'd6428, 25'd4761, 25'd1309, -25'd6666, -25'd5357}, '{25'd5476, -25'd119, 25'd12499, -25'd6666, -25'd4642, -25'd357, -25'd7975, 25'd1786, 25'd8332}, '{-25'd2619, 25'd12499, -25'd6666, -25'd833, 25'd13570, 25'd8570, 25'd1666, -25'd5118, 25'd4285}, '{25'd5595, -25'd4999, 25'd9761, -25'd2381, 25'd9047, -25'd4285, 25'd2976, 25'd6309, 25'd5118}, '{25'd3333, 25'd8332, -25'd7856, -25'd5952, -25'd2143, -25'd8332, 25'd5833, 25'd3214, 25'd7499}}},
    '{'{'{25'd15695, 25'd3488, -25'd698, 25'd1744, -25'd698, 25'd9591, -25'd6627, 25'd7150, -25'd2093}, '{-25'd2093, 25'd10114, 25'd11858, -25'd2790, 25'd3662, -25'd5232, -25'd5232, -25'd872, -25'd698}, '{-25'd1569, 25'd8370, -25'd8196, -25'd2616, 25'd10463, -25'd10986, -25'd4185, -25'd7847, 25'd11858}, '{-25'd2093, 25'd12730, 25'd3488, -25'd3139, 25'd12207, -25'd8545, 25'd6801, 25'd1395, -25'd872}, '{25'd5232, 25'd11335, 25'd1569, -25'd1046, 25'd5580, 25'd6452, 25'd5406, 25'd13602, 25'd5057}, '{-25'd523, 25'd349, -25'd2616, -25'd10637, -25'd4011, 25'd12032, 25'd4708, -25'd523, 25'd6103}, '{-25'd3139, -25'd4708, -25'd3488, 25'd5232, 25'd4185, 25'd11684, -25'd4185, -25'd9591, -25'd5232}, '{-25'd4883, -25'd12207, -25'd13428, -25'd2616, 25'd1569, -25'd14997, -25'd12556, -25'd9242, -25'd1221}, '{-25'd10114, -25'd3662, -25'd3662, -25'd20577, 25'd2616, -25'd8545, -25'd4011, -25'd2267, -25'd11684}}, '{'{-25'd8022, 25'd10289, 25'd3662, -25'd14299, -25'd8719, -25'd8370, 25'd174, -25'd14299, 25'd5057}, '{-25'd7847, -25'd4883, 25'd8196, -25'd1744, -25'd7324, -25'd14997, -25'd12730, 25'd1046, -25'd15695}, '{-25'd9765, 25'd6278, 25'd8196, 25'd3313, -25'd10289, -25'd3313, -25'd2616, -25'd1395, -25'd11684}, '{25'd12556, 25'd2790, -25'd174, -25'd11161, 25'd349, -25'd4360, -25'd9940, -25'd3662, 25'd5755}, '{-25'd1744, -25'd3662, -25'd9068, -25'd2093, -25'd1221, -25'd7498, 25'd2441, -25'd2790, -25'd7847}, '{-25'd2093, 25'd5755, -25'd8545, 25'd3139, 25'd5406, -25'd2616, -25'd7498, 25'd1395, 25'd5929}, '{25'd5580, -25'd8719, -25'd5232, -25'd8894, 25'd6278, 25'd2093, 25'd872, 25'd9591, 25'd698}, '{-25'd21100, -25'd15171, 25'd698, 25'd1744, -25'd2267, 25'd13602, 25'd1395, 25'd7150, -25'd2965}, '{-25'd15346, -25'd6103, 25'd11684, 25'd7150, 25'd10986, 25'd872, -25'd5057, -25'd7498, 25'd7847}}, '{'{25'd3662, -25'd6103, 25'd7847, -25'd2267, 25'd9417, 25'd3836, 25'd9765, 25'd8894, -25'd2965}, '{25'd10114, -25'd698, -25'd3836, -25'd13602, 25'd4011, 25'd3488, 25'd6801, 25'd1744, 25'd4360}, '{-25'd5406, 25'd8894, 25'd3139, 25'd5232, -25'd6627, 25'd2790, -25'd2965, 25'd5057, -25'd6627}, '{-25'd5057, 25'd1569, 25'd9417, -25'd8894, 25'd4360, -25'd5929, 25'd1744, 25'd1569, 25'd6801}, '{25'd5232, -25'd4883, -25'd523, -25'd10289, 25'd4185, 25'd9068, -25'd7324, -25'd7150, 25'd6103}, '{25'd9417, 25'd7324, -25'd3836, -25'd14823, -25'd5057, 25'd3662, 25'd9417, -25'd3662, -25'd13951}, '{-25'd7324, -25'd14299, -25'd3139, 25'd5057, 25'd5929, 25'd9940, 25'd3836, 25'd5406, 25'd4883}, '{-25'd12381, -25'd21449, -25'd17613, -25'd22147, -25'd2790, -25'd3313, -25'd523, -25'd8545, 25'd4883}, '{-25'd1046, -25'd13776, -25'd16043, -25'd21449, 25'd9068, 25'd12032, 25'd5406, -25'd5057, -25'd4360}}},
    '{'{'{-25'd4743, -25'd6838, -25'd8824, 25'd1544, 25'd6507, -25'd8713, -25'd4412, 25'd6728, 25'd221}, '{-25'd1434, 25'd10588, 25'd6507, 25'd3640, 25'd9044, 25'd4632, 25'd6397, -25'd6507, -25'd9485}, '{-25'd441, 25'd1875, -25'd882, 25'd10037, -25'd1544, 25'd8934, 25'd9816, 25'd1103, 25'd14007}, '{-25'd441, 25'd8382, 25'd11250, -25'd7941, -25'd5074, 25'd8713, -25'd2206, -25'd993, 25'd5846}, '{-25'd7610, -25'd2537, -25'd11912, 25'd5515, 25'd1324, 25'd11360, -25'd3199, -25'd3971, 25'd2096}, '{-25'd6066, 25'd8713, -25'd4081, -25'd9044, 25'd1434, -25'd7721, 25'd10478, 25'd5184, -25'd7059}, '{-25'd1324, 25'd9375, 25'd5294, 25'd110, 25'd2757, 25'd1985, 25'd4632, 25'd9816, -25'd1324}, '{-25'd6066, -25'd10478, -25'd4632, -25'd1985, -25'd7169, -25'd10368, 25'd110, 25'd8162, -25'd11250}, '{-25'd10147, 25'd6838, -25'd4081, -25'd2868, -25'd8162, -25'd10368, 25'd1324, 25'd4522, -25'd7610}}, '{'{25'd9706, -25'd551, 25'd9485, 25'd11581, 25'd8824, 25'd11912, -25'd772, 25'd9926, 25'd4081}, '{25'd8493, -25'd2096, -25'd3750, -25'd10147, 25'd11029, -25'd5515, 25'd11250, -25'd9265, -25'd3199}, '{-25'd4081, -25'd5074, 25'd8272, 25'd3529, 25'd3419, -25'd2096, -25'd8272, 25'd9375, -25'd4743}, '{25'd1103, 25'd1324, -25'd12463, 25'd3419, 25'd11801, -25'd1213, -25'd10368, 25'd8713, -25'd662}, '{25'd441, 25'd4853, 25'd5184, -25'd4081, -25'd1544, 25'd1985, 25'd7279, -25'd2978, 25'd11140}, '{-25'd1875, -25'd5184, -25'd5294, 25'd5074, 25'd772, 25'd882, 25'd10368, 25'd1544, 25'd5735}, '{-25'd5074, 25'd9375, 25'd3640, -25'd11360, -25'd11581, -25'd9816, 25'd10478, 25'd2426, 25'd1765}, '{25'd8272, -25'd13015, -25'd8382, -25'd4522, 25'd10257, -25'd2868, 25'd1765, 25'd5294, -25'd3419}, '{25'd4191, -25'd9044, -25'd2537, 25'd10257, -25'd6507, -25'd4632, -25'd11691, -25'd7941, 25'd3860}}, '{'{25'd4632, 25'd9044, 25'd3971, -25'd2316, 25'd7279, -25'd4522, -25'd6838, 25'd11250, 25'd12573}, '{25'd8051, 25'd7169, 25'd3529, -25'd10698, 25'd10809, -25'd6397, -25'd1765, -25'd882, 25'd7390}, '{-25'd11912, 25'd11029, 25'd7279, -25'd8603, 25'd1875, -25'd2537, 25'd10147, 25'd11360, -25'd4191}, '{25'd4081, 25'd11360, 25'd11029, 25'd3750, 25'd10698, -25'd7279, 25'd7610, 25'd7169, -25'd1875}, '{25'd2426, 25'd662, -25'd3309, 25'd2757, -25'd1213, -25'd772, 25'd5846, -25'd3309, -25'd7500}, '{25'd8162, 25'd9044, -25'd7500, -25'd5846, -25'd1544, 25'd6507, -25'd3640, -25'd6066, -25'd10478}, '{25'd8382, -25'd7059, -25'd5956, -25'd6287, -25'd6618, -25'd8824, -25'd4301, -25'd11029, 25'd10809}, '{-25'd11801, -25'd10037, -25'd8162, 25'd7721, 25'd1654, 25'd1765, -25'd10919, 25'd5625, 25'd1434}, '{-25'd3199, 25'd4191, -25'd5074, 25'd551, -25'd4522, 25'd6507, 25'd6176, -25'd3640, -25'd11581}}},
    '{'{'{-25'd4072, 25'd10502, 25'd8573, 25'd8787, 25'd11788, 25'd7930, -25'd7501, 25'd4394, 25'd3536}, '{-25'd1286, -25'd11788, 25'd4072, 25'd8251, 25'd8358, 25'd9644, -25'd3429, 25'd6108, 25'd11145}, '{-25'd107, 25'd1286, 25'd2358, 25'd9644, 25'd6430, -25'd1393, -25'd7180, 25'd4501, -25'd2893}, '{-25'd5358, 25'd3858, -25'd6537, -25'd5358, -25'd4072, -25'd10073, -25'd3429, -25'd8358, 25'd1607}, '{-25'd3322, -25'd214, -25'd7394, 25'd9859, 25'd10073, -25'd9966, -25'd5679, 25'd857, 25'd8037}, '{-25'd6644, -25'd10287, 25'd2036, 25'd4929, 25'd8894, 25'd4286, -25'd2679, 25'd7180, 25'd2143}, '{25'd10502, 25'd7501, -25'd2679, -25'd7715, -25'd964, -25'd4072, -25'd5358, 25'd5465, -25'd11252}, '{-25'd8787, 25'd1286, 25'd7823, -25'd8466, 25'd7823, 25'd214, 25'd1179, -25'd1822, -25'd321}, '{25'd3858, 25'd5465, 25'd1607, -25'd1607, -25'd10287, 25'd5358, -25'd4929, -25'd4822, -25'd4608}}, '{'{-25'd11037, -25'd1607, -25'd10502, -25'd9216, 25'd4929, 25'd6644, -25'd10073, 25'd8251, 25'd9430}, '{-25'd6858, -25'd9537, 25'd7501, -25'd10287, -25'd3643, -25'd4822, -25'd6215, -25'd1072, -25'd9751}, '{-25'd12002, -25'd750, -25'd11466, 25'd9323, 25'd4179, -25'd4715, -25'd11466, 25'd10287, -25'd4394}, '{-25'd1715, -25'd8573, -25'd3108, 25'd9001, -25'd6001, -25'd1286, 25'd2036, 25'd750, 25'd10716}, '{-25'd964, 25'd1607, 25'd10930, -25'd8358, -25'd10502, 25'd1179, 25'd8251, -25'd5679, -25'd1715}, '{-25'd10930, -25'd12216, 25'd7180, 25'd12430, 25'd429, 25'd3000, 25'd8894, 25'd10073, -25'd4179}, '{-25'd10287, 25'd1500, 25'd7073, 25'd4501, 25'd9216, -25'd4072, -25'd10716, -25'd1179, -25'd3643}, '{-25'd3000, -25'd1072, -25'd11680, 25'd9644, 25'd7180, 25'd0, 25'd9216, -25'd1286, 25'd8251}, '{-25'd9751, -25'd1715, 25'd8251, 25'd1179, -25'd8680, 25'd1715, -25'd10930, -25'd2786, -25'd3215}}, '{'{-25'd2465, -25'd7823, -25'd9323, -25'd1286, -25'd8894, 25'd5036, -25'd750, -25'd11252, -25'd3000}, '{-25'd9537, -25'd6430, 25'd2143, -25'd9537, 25'd7823, -25'd4929, -25'd429, 25'd9751, 25'd7180}, '{-25'd10394, -25'd7394, -25'd3215, 25'd8144, -25'd2679, 25'd1822, 25'd9323, -25'd3429, -25'd11359}, '{-25'd1500, -25'd13716, -25'd5894, 25'd0, -25'd9216, 25'd1715, -25'd1607, 25'd7394, -25'd964}, '{25'd4608, -25'd6858, 25'd857, 25'd7180, 25'd107, 25'd5679, -25'd5465, 25'd8680, 25'd5144}, '{-25'd3322, 25'd7394, 25'd4608, 25'd10823, -25'd5144, 25'd2572, -25'd3643, 25'd3858, 25'd3215}, '{-25'd8251, -25'd10609, 25'd7608, 25'd8680, 25'd10287, -25'd4286, -25'd4929, 25'd5894, 25'd11037}, '{25'd4929, -25'd4929, -25'd8144, -25'd5251, -25'd11145, 25'd9751, -25'd9323, -25'd8573, 25'd1179}, '{-25'd7823, 25'd4286, 25'd9323, 25'd2465, 25'd1929, 25'd429, 25'd9859, 25'd6965, -25'd3643}}},
    '{'{'{-25'd11044, 25'd7233, 25'd7233, -25'd7819, -25'd6158, -25'd4789, -25'd684, 25'd6548, 25'd6646}, '{-25'd3519, 25'd4594, 25'd10751, -25'd3616, 25'd1271, 25'd6842, 25'd5669, -25'd9774, -25'd1759}, '{-25'd2541, 25'd11044, -25'd9676, -25'd11044, -25'd3812, -25'd6548, -25'd4496, -25'd3030, -25'd3323}, '{25'd4789, 25'd1759, 25'd391, 25'd3128, 25'd489, -25'd6842, -25'd9774, -25'd8796, -25'd6451}, '{-25'd4594, 25'd11240, 25'd4007, -25'd5669, -25'd489, -25'd10653, -25'd1955, -25'd8406, 25'd6255}, '{25'd8796, 25'd8894, -25'd391, 25'd9578, 25'd2443, 25'd3714, -25'd2248, 25'd4985, -25'd7330}, '{-25'd7721, 25'd9872, -25'd5278, -25'd8308, -25'd2346, 25'd5180, -25'd6451, -25'd1564, 25'd6060}, '{-25'd4594, -25'd10556, 25'd195, 25'd293, -25'd4594, -25'd684, -25'd3421, 25'd7819, 25'd8308}, '{25'd293, 25'd1564, 25'd10067, 25'd11044, -25'd4300, 25'd9481, -25'd8992, 25'd11435, -25'd9676}}, '{'{25'd4496, 25'd11338, 25'd1368, -25'd3030, -25'd3421, -25'd9481, -25'd1368, -25'd98, 25'd6353}, '{-25'd5082, -25'd7819, 25'd3616, 25'd3812, 25'd2834, 25'd11826, 25'd4887, 25'd9578, 25'd9774}, '{-25'd3812, 25'd8015, 25'd6548, -25'd2639, 25'd10653, 25'd10751, 25'd7330, 25'd11533, -25'd1368}, '{-25'd6451, -25'd10263, -25'd10360, 25'd6939, -25'd6842, 25'd10458, -25'd2639, -25'd4398, 25'd5669}, '{-25'd4887, 25'd4007, -25'd4496, -25'd8601, 25'd11729, -25'd6744, 25'd7135, -25'd782, 25'd977}, '{25'd9774, -25'd11338, -25'd10458, 25'd5669, 25'd1368, -25'd6060, 25'd10556, 25'd7819, -25'd6842}, '{25'd1857, -25'd11142, -25'd6451, -25'd4007, -25'd4887, 25'd6939, 25'd1759, 25'd5571, 25'd880}, '{25'd5473, -25'd3030, -25'd1564, 25'd1368, 25'd4691, -25'd8992, 25'd9187, 25'd2834, 25'd3323}, '{25'd3225, -25'd4594, -25'd6744, -25'd10067, 25'd12217, -25'd8796, 25'd4203, -25'd4105, 25'd6158}}, '{'{-25'd4691, 25'd5376, 25'd5669, 25'd8601, 25'd2541, -25'd4985, -25'd10458, -25'd11044, -25'd4887}, '{25'd5767, 25'd11240, 25'd7819, -25'd8308, 25'd4007, -25'd9285, -25'd2737, 25'd8699, 25'd6451}, '{-25'd5571, 25'd12413, -25'd11631, -25'd8992, -25'd10556, 25'd10849, 25'd7917, -25'd3812, 25'd4007}, '{-25'd8015, 25'd11631, -25'd391, 25'd0, 25'd7330, 25'd8112, -25'd4300, 25'd2053, -25'd12120}, '{-25'd5864, 25'd2248, 25'd11142, 25'd2834, 25'd9187, 25'd7819, 25'd1466, -25'd8699, -25'd1955}, '{25'd2737, -25'd3128, 25'd7526, -25'd4887, -25'd9872, 25'd6353, 25'd2443, -25'd2834, 25'd195}, '{-25'd7721, 25'd1955, 25'd11142, -25'd6353, 25'd6744, 25'd3519, -25'd782, 25'd11142, 25'd4789}, '{25'd4594, 25'd1564, 25'd11338, -25'd8406, 25'd3519, 25'd1173, 25'd7428, 25'd9969, -25'd6158}, '{-25'd10165, -25'd5669, 25'd10458, -25'd11142, -25'd6646, 25'd1173, 25'd9481, -25'd10653, 25'd3128}}},
    '{'{'{-25'd1559, 25'd10812, -25'd7797, 25'd1559, 25'd9668, 25'd1871, -25'd6342, -25'd8941, 25'd6134}, '{-25'd6861, 25'd11332, 25'd10604, -25'd312, 25'd7485, 25'd6654, 25'd5614, 25'd8109, -25'd12060}, '{25'd7069, 25'd8941, -25'd8005, 25'd6342, 25'd3431, -25'd5406, 25'd9980, -25'd624, -25'd4158}, '{-25'd3223, 25'd3223, -25'd10916, -25'd12268, -25'd11852, 25'd728, 25'd7069, 25'd2391, -25'd11332}, '{-25'd4470, 25'd312, 25'd7069, 25'd10604, 25'd1352, 25'd8837, -25'd13203, -25'd8317, 25'd1455}, '{-25'd10604, -25'd6965, -25'd9668, 25'd3639, 25'd832, 25'd5926, -25'd6654, 25'd6134, 25'd2183}, '{25'd6654, -25'd9149, 25'd10604, 25'd4574, -25'd8421, 25'd4262, -25'd11124, 25'd5718, -25'd12164}, '{-25'd9772, 25'd8005, -25'd1559, -25'd10708, -25'd3223, -25'd7381, -25'd12371, -25'd7173, 25'd1975}, '{-25'd9461, 25'd3743, 25'd6342, -25'd10916, -25'd7173, 25'd2911, 25'd9876, -25'd11748, -25'd1871}}, '{'{-25'd3743, -25'd9149, -25'd3327, 25'd8629, 25'd4678, -25'd8109, 25'd11124, -25'd7485, -25'd936}, '{25'd4886, 25'd8525, 25'd11748, 25'd5406, 25'd8317, 25'd4262, 25'd10188, 25'd5302, 25'd3535}, '{25'd9772, -25'd9357, -25'd3431, 25'd3951, -25'd9357, -25'd416, -25'd416, -25'd1248, 25'd11228}, '{-25'd7277, -25'd10916, 25'd10916, 25'd9668, 25'd9149, 25'd4678, 25'd11020, 25'd4678, -25'd1248}, '{25'd6238, 25'd6030, 25'd2807, -25'd6550, -25'd2599, -25'd8421, 25'd6446, 25'd1248, -25'd6134}, '{-25'd9253, -25'd8005, 25'd4055, -25'd8837, -25'd6965, -25'd1767, -25'd3847, -25'd12060, 25'd10396}, '{25'd1871, -25'd9045, 25'd5926, 25'd6654, 25'd4158, -25'd4574, -25'd4574, -25'd6238, 25'd5718}, '{25'd8213, 25'd104, -25'd1663, -25'd624, -25'd6446, -25'd9980, -25'd8837, -25'd12268, -25'd9045}, '{-25'd8213, -25'd7173, 25'd3639, 25'd1559, 25'd9668, -25'd832, -25'd832, -25'd12060, -25'd4678}}, '{'{25'd10708, 25'd6550, 25'd11228, 25'd1248, -25'd7901, 25'd10188, -25'd832, -25'd8629, 25'd9045}, '{25'd4782, 25'd8317, 25'd11124, 25'd5406, -25'd6550, -25'd3535, 25'd12787, 25'd11436, 25'd12164}, '{25'd10396, 25'd4886, -25'd10604, 25'd3119, 25'd10916, 25'd1767, 25'd208, 25'd5614, -25'd7797}, '{-25'd7381, 25'd4678, 25'd5094, 25'd5822, 25'd6965, 25'd7485, -25'd6238, 25'd7069, -25'd8109}, '{25'd9772, -25'd1767, 25'd8421, 25'd2807, -25'd8109, 25'd8317, -25'd9149, 25'd3639, 25'd5510}, '{25'd6550, -25'd11332, 25'd12060, 25'd7693, -25'd9045, 25'd5406, 25'd12164, 25'd6134, 25'd5094}, '{-25'd10708, 25'd9668, 25'd11020, 25'd11956, -25'd6965, 25'd8213, 25'd5614, 25'd5926, 25'd2495}, '{-25'd6654, -25'd6861, -25'd3431, 25'd624, 25'd6758, 25'd2079, -25'd6654, -25'd5614, -25'd8837}, '{25'd4990, 25'd10500, -25'd2183, -25'd3015, 25'd2183, -25'd10084, 25'd7901, 25'd8317, 25'd11748}}},
    '{'{'{25'd5847, -25'd5630, -25'd1732, -25'd4981, -25'd3790, 25'd4223, -25'd8120, -25'd2165, 25'd3465}, '{-25'd2599, -25'd2057, -25'd9853, -25'd1624, 25'd3898, 25'd0, 25'd5305, 25'd11910, 25'd12560}, '{25'd1949, -25'd217, -25'd10069, 25'd11802, -25'd9203, 25'd11369, -25'd2707, -25'd2707, 25'd8229}, '{25'd0, 25'd3356, 25'd6605, 25'd2923, -25'd10719, -25'd10611, -25'd9853, -25'd6605, -25'd325}, '{25'd11585, -25'd9095, 25'd8553, -25'd1083, -25'd10286, -25'd433, -25'd5522, -25'd1516, 25'd11260}, '{-25'd7038, -25'd5305, 25'd7904, 25'd3573, 25'd9744, -25'd2057, 25'd7904, -25'd5305, -25'd9095}, '{-25'd1841, -25'd4547, 25'd4547, -25'd8012, -25'd4114, -25'd2490, 25'd11477, 25'd4114, -25'd7796}, '{25'd11369, 25'd8337, 25'd3356, 25'd4547, -25'd1949, 25'd12884, 25'd7038, -25'd6063, -25'd7904}, '{25'd9203, 25'd2382, -25'd4223, -25'd4223, -25'd8012, 25'd2490, -25'd3573, -25'd9420, 25'd2923}}, '{'{-25'd4439, 25'd9636, 25'd5197, -25'd2707, -25'd4006, -25'd3681, -25'd7904, 25'd1408, -25'd2057}, '{-25'd5847, 25'd7363, 25'd5197, 25'd0, 25'd7904, -25'd8987, 25'd10611, 25'd10827, -25'd8662}, '{25'd5089, 25'd9528, -25'd1732, -25'd3356, 25'd4331, 25'd3898, -25'd9744, 25'd3898, -25'd4656}, '{25'd4331, 25'd3681, -25'd2057, 25'd3248, -25'd8120, -25'd866, 25'd7471, -25'd3573, 25'd8012}, '{25'd8770, 25'd325, -25'd541, -25'd2599, -25'd5630, -25'd6605, 25'd0, 25'd4547, 25'd8770}, '{-25'd3790, -25'd7904, -25'd4764, -25'd2707, -25'd3898, -25'd5197, -25'd2490, -25'd3032, 25'd12126}, '{-25'd5847, -25'd4331, -25'd11044, 25'd9528, -25'd4331, -25'd8445, 25'd7579, -25'd4331, -25'd10935}, '{25'd7146, -25'd4547, 25'd7904, -25'd325, -25'd9744, 25'd10069, 25'd10611, -25'd2923, 25'd1516}, '{-25'd4981, 25'd3356, 25'd8229, 25'd9095, 25'd12126, -25'd6605, -25'd1516, -25'd974, -25'd3681}}, '{'{-25'd8553, 25'd4981, 25'd8229, 25'd3898, 25'd8987, 25'd11260, 25'd12343, 25'd13426, 25'd9528}, '{25'd6388, 25'd8662, 25'd974, 25'd1732, 25'd6929, -25'd7363, 25'd9636, -25'd6063, 25'd2274}, '{25'd7363, -25'd3140, 25'd7363, 25'd4764, 25'd6605, 25'd12884, 25'd5414, -25'd4114, 25'd13751}, '{25'd2599, 25'd4764, 25'd541, 25'd11152, -25'd9636, 25'd4547, -25'd5522, 25'd10178, 25'd1299}, '{25'd7254, 25'd2815, 25'd9311, -25'd541, -25'd7146, 25'd4656, 25'd4872, 25'd6605, -25'd6280}, '{25'd7363, -25'd3790, -25'd8229, -25'd9311, 25'd217, 25'd11585, 25'd6605, -25'd5414, 25'd758}, '{25'd6713, -25'd3573, -25'd9311, -25'd10178, 25'd1732, -25'd3356, -25'd2490, 25'd8229, -25'd2490}, '{25'd4547, -25'd2382, 25'd1408, 25'd9420, 25'd4006, -25'd7038, 25'd5197, -25'd8012, 25'd5630}, '{-25'd1083, 25'd9528, 25'd11044, 25'd7904, -25'd4439, 25'd3356, -25'd7146, -25'd8662, -25'd3681}}},
    '{'{'{-25'd8351, 25'd6236, 25'd0, -25'd1448, 25'd1448, 25'd668, 25'd8129, -25'd2227, -25'd10578}, '{25'd8240, 25'd4899, -25'd6347, -25'd11469, -25'd1114, -25'd12360, 25'd334, 25'd2784, -25'd4454}, '{25'd7461, 25'd1336, 25'd6458, 25'd1114, -25'd1893, 25'd8351, -25'd3675, 25'd223, 25'd6458}, '{-25'd4009, 25'd8017, 25'd8908, -25'd1448, 25'd1782, -25'd5122, 25'd10244, -25'd8908, -25'd11692}, '{25'd6236, 25'd6124, -25'd7349, -25'd5011, -25'd9576, -25'd11358, 25'd7238, -25'd8797, -25'd4231}, '{-25'd6681, -25'd668, 25'd8129, -25'd12471, -25'd2227, -25'd6570, 25'd8685, 25'd4454, -25'd5790}, '{25'd10356, -25'd3452, -25'd1893, 25'd3229, -25'd9354, 25'd2338, -25'd6124, -25'd3675, 25'd4343}, '{-25'd11469, -25'd9242, 25'd8240, -25'd9354, 25'd10356, -25'd7906, -25'd6792, -25'd9688, 25'd6792}, '{25'd8463, -25'd8797, -25'd1893, -25'd5456, 25'd5345, 25'd7238, -25'd8574, 25'd2116, 25'd2338}}, '{'{25'd5568, -25'd7906, 25'd1002, 25'd5790, -25'd3229, -25'd1114, -25'd14253, -25'd2561, 25'd5122}, '{25'd6570, 25'd668, -25'd13474, -25'd5902, -25'd14253, -25'd13251, 25'd5122, 25'd4343, -25'd11581}, '{-25'd9799, -25'd2450, -25'd3897, -25'd9354, -25'd111, 25'd6792, -25'd10244, -25'd10022, -25'd8685}, '{-25'd5790, 25'd6681, -25'd5568, 25'd2227, -25'd11247, -25'd6792, 25'd7461, -25'd2561, -25'd8685}, '{-25'd5456, 25'd5234, -25'd10912, 25'd2450, -25'd7572, 25'd4231, -25'd7795, -25'd12249, -25'd13251}, '{-25'd11469, -25'd6681, 25'd5011, 25'd1782, -25'd8351, -25'd12137, -25'd5234, -25'd11135, -25'd11135}, '{-25'd8351, -25'd1893, 25'd1114, -25'd7015, 25'd1893, 25'd1336, 25'd4231, 25'd1670, -25'd2895}, '{25'd2672, -25'd13808, 25'd7349, 25'd668, -25'd9354, -25'd11803, 25'd7906, -25'd8017, -25'd10912}, '{-25'd9131, 25'd8351, -25'd12694, -25'd4565, 25'd5011, -25'd8574, -25'd1893, 25'd8351, -25'd1336}}, '{'{25'd3229, -25'd5345, 25'd7683, -25'd6792, 25'd4565, 25'd12137, 25'd3563, 25'd11581, 25'd4454}, '{25'd13696, 25'd12360, 25'd8017, -25'd8574, 25'd4899, 25'd10912, -25'd2116, -25'd1670, -25'd8240}, '{25'd12360, -25'd9242, 25'd1114, -25'd7015, -25'd10578, 25'd3452, 25'd3341, -25'd9465, 25'd9688}, '{25'd9688, 25'd7015, 25'd10467, 25'd11915, 25'd4788, -25'd1225, -25'd7906, 25'd8129, 25'd6681}, '{25'd7349, -25'd10022, -25'd6904, 25'd3675, -25'd9354, 25'd9354, -25'd6570, -25'd5456, 25'd1336}, '{-25'd4565, -25'd7349, -25'd11135, 25'd9465, -25'd9354, -25'd223, -25'd9576, 25'd779, 25'd4788}, '{25'd10022, 25'd6347, 25'd2450, -25'd6681, -25'd1114, -25'd4120, -25'd5790, -25'd2895, 25'd13028}, '{-25'd891, 25'd5568, -25'd9354, -25'd4231, 25'd3897, 25'd12360, -25'd334, 25'd4343, 25'd6013}, '{25'd0, 25'd12805, -25'd3675, -25'd668, -25'd5790, 25'd4454, 25'd0, -25'd6792, -25'd1225}}},
    '{'{'{25'd106, 25'd9667, -25'd9348, 25'd6480, 25'd9454, 25'd5949, -25'd3187, 25'd8073, 25'd3824}, '{-25'd4143, 25'd13066, 25'd7967, -25'd7011, 25'd7861, -25'd637, -25'd6799, 25'd744, 25'd637}, '{25'd7224, 25'd6055, 25'd5630, 25'd10304, 25'd3399, 25'd7117, 25'd10198, -25'd956, -25'd2018}, '{25'd8498, -25'd1593, 25'd8605, -25'd9561, -25'd4568, -25'd8817, -25'd6480, -25'd531, -25'd10198}, '{-25'd3187, 25'd3081, 25'd7117, 25'd11791, 25'd3824, 25'd10092, -25'd4462, 25'd1381, 25'd7542}, '{-25'd5311, 25'd10729, 25'd9879, 25'd9986, 25'd5736, -25'd8392, 25'd13066, -25'd1806, -25'd3612}, '{25'd3824, 25'd12110, 25'd5630, 25'd5205, -25'd7542, -25'd3506, 25'd10729, 25'd2125, 25'd10729}, '{-25'd425, -25'd3187, 25'd11048, 25'd744, 25'd8286, 25'd1169, -25'd5205, -25'd2549, 25'd5524}, '{25'd3612, 25'd4037, 25'd8817, 25'd8392, 25'd11154, -25'd744, -25'd4249, -25'd4462, 25'd12323}}, '{'{-25'd12429, -25'd13279, 25'd3824, 25'd850, 25'd9242, -25'd13491, -25'd7755, 25'd1275, -25'd4355}, '{-25'd744, -25'd7861, 25'd3081, 25'd9348, -25'd4887, 25'd3612, -25'd6480, -25'd9879, -25'd425}, '{-25'd3187, -25'd1169, -25'd10410, 25'd8392, -25'd4568, 25'd2125, -25'd6799, -25'd11260, -25'd4993}, '{-25'd9242, 25'd5099, 25'd2868, -25'd6374, -25'd9029, 25'd1806, 25'd5949, -25'd9348, 25'd5418}, '{25'd1593, 25'd744, -25'd1806, -25'd6267, -25'd1912, -25'd7330, -25'd9136, -25'd1806, 25'd8073}, '{25'd5418, -25'd8286, 25'd4249, 25'd8073, -25'd2018, 25'd956, -25'd10942, 25'd212, -25'd7436}, '{25'd8392, 25'd8286, 25'd2337, 25'd9667, 25'd8073, 25'd5736, 25'd11473, 25'd9561, -25'd956}, '{-25'd3718, 25'd9773, -25'd1275, 25'd4462, -25'd637, 25'd3824, -25'd6374, -25'd212, 25'd8180}, '{25'd1487, -25'd2337, -25'd3718, 25'd2337, -25'd12110, 25'd2974, -25'd9773, 25'd10623, -25'd11048}}, '{'{-25'd6055, -25'd744, -25'd5099, 25'd212, 25'd6905, 25'd6799, 25'd12110, 25'd5524, -25'd3506}, '{-25'd3399, 25'd1593, 25'd10410, -25'd8286, -25'd7542, 25'd12747, -25'd8605, -25'd1700, -25'd8286}, '{-25'd10835, -25'd2868, 25'd5205, 25'd10623, -25'd2656, -25'd10410, 25'd1912, -25'd2868, -25'd5949}, '{-25'd212, -25'd7861, -25'd2762, -25'd4355, 25'd5736, -25'd744, -25'd9986, 25'd5843, -25'd5736}, '{25'd2231, 25'd9561, 25'd4568, 25'd4462, -25'd11048, 25'd11048, 25'd1275, 25'd9561, -25'd7224}, '{25'd3824, -25'd1275, -25'd10942, 25'd8817, -25'd1381, -25'd1381, -25'd8605, -25'd4568, -25'd9773}, '{-25'd9029, 25'd11473, 25'd1806, 25'd7967, -25'd9667, 25'd4462, -25'd3399, 25'd3718, -25'd1062}, '{25'd1169, -25'd4568, -25'd12110, -25'd8711, -25'd5630, -25'd5418, -25'd4887, -25'd12004, 25'd8711}, '{25'd5311, 25'd3930, -25'd12004, 25'd8498, -25'd5099, 25'd1806, -25'd12004, 25'd10835, 25'd9773}}},
    '{'{'{25'd3691, -25'd13262, 25'd2051, 25'd6836, 25'd11621, 25'd3418, 25'd12031, 25'd2051, 25'd8613}, '{25'd1914, -25'd2871, -25'd820, 25'd9980, 25'd9023, -25'd8203, 25'd547, -25'd1094, 25'd2324}, '{25'd10117, -25'd10117, -25'd9297, 25'd9844, 25'd4922, 25'd6562, -25'd6016, 25'd7383, 25'd11348}, '{25'd1504, 25'd5742, 25'd7656, 25'd6973, 25'd6426, 25'd12851, 25'd3008, -25'd1914, 25'd957}, '{25'd6016, -25'd8887, 25'd7246, 25'd7109, 25'd6836, -25'd8750, -25'd4238, 25'd14082, -25'd4922}, '{25'd9844, -25'd9160, -25'd547, -25'd10117, 25'd820, -25'd1641, -25'd5605, -25'd8476, 25'd5059}, '{25'd9023, -25'd3555, -25'd5195, -25'd5469, 25'd13398, -25'd8340, -25'd6152, 25'd12441, 25'd1641}, '{-25'd9707, 25'd12578, -25'd3965, 25'd9844, -25'd9844, 25'd9160, 25'd5879, -25'd7656, -25'd8066}, '{-25'd9980, 25'd4512, -25'd5605, 25'd3828, 25'd2187, 25'd11211, -25'd8340, 25'd273, -25'd9297}}, '{'{-25'd2324, 25'd5332, -25'd2461, 25'd5332, 25'd3008, -25'd11894, -25'd3281, 25'd547, -25'd7383}, '{-25'd11074, -25'd2187, -25'd15176, -25'd14355, -25'd10254, -25'd13945, -25'd6152, -25'd4238, -25'd9707}, '{-25'd6562, 25'd5742, -25'd15996, 25'd7656, 25'd1777, -25'd5879, 25'd8066, -25'd9844, -25'd9844}, '{-25'd5879, -25'd12168, -25'd17500, -25'd12715, -25'd14492, -25'd12305, 25'd820, -25'd11758, -25'd7930}, '{-25'd10527, -25'd957, 25'd4512, -25'd2734, 25'd8476, 25'd3555, 25'd1641, 25'd0, -25'd12578}, '{-25'd14629, 25'd5332, -25'd12851, -25'd410, -25'd8750, -25'd3145, 25'd1367, 25'd9434, 25'd4922}, '{-25'd9160, -25'd12168, -25'd10117, 25'd7246, 25'd820, -25'd8340, 25'd1230, -25'd4375, -25'd5469}, '{-25'd5059, -25'd12715, -25'd13398, 25'd8203, -25'd2324, 25'd7930, 25'd3418, -25'd2461, -25'd5059}, '{-25'd2324, -25'd3555, -25'd8203, 25'd8887, 25'd9160, -25'd4785, 25'd9297, 25'd410, -25'd2461}}, '{'{-25'd4375, -25'd10254, -25'd8750, -25'd3418, 25'd1230, 25'd4102, -25'd8203, 25'd11211, 25'd6836}, '{25'd8750, 25'd410, 25'd11621, 25'd6016, -25'd8066, 25'd13398, 25'd6562, 25'd8066, -25'd820}, '{-25'd1777, -25'd10391, -25'd9023, -25'd9297, -25'd1641, 25'd6562, -25'd7793, 25'd12441, 25'd3008}, '{25'd9297, 25'd5742, 25'd2461, 25'd9844, -25'd9434, 25'd7656, 25'd12031, 25'd8750, -25'd5059}, '{-25'd2324, -25'd7930, -25'd7656, 25'd13808, -25'd6699, -25'd273, 25'd12441, -25'd2051, -25'd1914}, '{25'd5605, -25'd5742, 25'd12031, 25'd5469, -25'd5332, 25'd7793, -25'd2324, 25'd4375, 25'd8887}, '{-25'd5879, -25'd6699, -25'd4922, 25'd14355, 25'd4375, 25'd10527, 25'd9570, 25'd9160, 25'd13398}, '{25'd7930, 25'd10117, -25'd3691, 25'd4375, -25'd2871, -25'd4785, 25'd9570, 25'd12031, 25'd6973}, '{25'd11894, -25'd5332, 25'd13808, 25'd14629, 25'd1777, -25'd8203, -25'd2871, -25'd7793, 25'd10801}}},
    '{'{'{25'd0, -25'd9262, -25'd9056, -25'd12555, 25'd8953, 25'd5043, -25'd5454, 25'd7204, 25'd2984}, '{25'd823, 25'd9777, 25'd8027, -25'd4528, -25'd12967, -25'd4631, 25'd3396, -25'd8542, -25'd5454}, '{-25'd10806, 25'd7101, 25'd8953, 25'd8233, -25'd12041, -25'd9571, 25'd7821, -25'd4940, -25'd3293}, '{25'd5557, -25'd11320, 25'd4117, 25'd2470, 25'd8130, -25'd4940, -25'd13173, 25'd3190, 25'd3602}, '{25'd5969, 25'd1235, -25'd12350, -25'd7101, 25'd8233, -25'd4631, 25'd3808, 25'd6895, 25'd4322}, '{-25'd8953, 25'd10085, 25'd617, -25'd2676, 25'd6586, 25'd823, -25'd2882, -25'd5660, 25'd1132}, '{25'd3190, 25'd7718, 25'd103, -25'd720, -25'd13070, -25'd1544, 25'd3602, 25'd10600, 25'd9983}, '{25'd5454, 25'd9983, -25'd11423, 25'd3087, -25'd4219, 25'd6895, 25'd7307, 25'd8748, -25'd2470}, '{25'd5660, -25'd10806, -25'd11835, -25'd5557, -25'd10291, 25'd6175, -25'd11938, -25'd6586, 25'd617}}, '{'{-25'd1338, -25'd7718, 25'd4631, 25'd4014, -25'd3190, 25'd2882, -25'd10497, 25'd103, 25'd617}, '{25'd3499, -25'd10806, 25'd6483, 25'd1955, 25'd5146, -25'd2676, -25'd5043, -25'd5763, -25'd103}, '{-25'd1544, -25'd12041, 25'd926, 25'd1852, -25'd1441, -25'd1132, 25'd7513, 25'd6278, -25'd11938}, '{-25'd11629, 25'd6483, -25'd5146, -25'd6278, 25'd1647, -25'd2882, 25'd9571, -25'd4425, -25'd2161}, '{-25'd4322, -25'd7616, -25'd12864, -25'd8233, 25'd309, 25'd10085, 25'd4528, 25'd7204, -25'd11423}, '{-25'd5351, 25'd2264, -25'd6998, -25'd10291, -25'd412, -25'd11012, 25'd926, 25'd1955, -25'd3602}, '{-25'd12041, -25'd10188, -25'd4837, 25'd8850, 25'd8542, -25'd10909, -25'd11732, 25'd9777, 25'd7513}, '{-25'd9262, 25'd823, -25'd1544, -25'd8542, -25'd12967, 25'd2676, -25'd5454, -25'd6278, -25'd4219}, '{-25'd1544, -25'd4014, 25'd6175, 25'd103, -25'd4425, 25'd6483, -25'd1029, -25'd11526, -25'd9365}}, '{'{-25'd5454, 25'd0, 25'd3499, 25'd2470, -25'd1338, 25'd3602, 25'd6483, 25'd4528, 25'd206}, '{-25'd1338, 25'd7616, -25'd1647, 25'd1544, 25'd1647, 25'd5351, 25'd103, 25'd3293, -25'd8027}, '{-25'd2264, -25'd6278, 25'd4528, -25'd6586, 25'd6278, -25'd8336, -25'd6998, -25'd3808, 25'd8645}, '{25'd6381, -25'd7616, -25'd9365, 25'd926, 25'd4734, -25'd1955, -25'd3911, 25'd926, 25'd9880}, '{25'd9262, -25'd2264, -25'd823, 25'd2779, -25'd5969, 25'd5043, 25'd5866, 25'd4528, 25'd6586}, '{-25'd11938, -25'd4219, -25'd823, -25'd10909, 25'd8336, -25'd1338, -25'd926, 25'd5969, 25'd5454}, '{-25'd7718, -25'd9365, 25'd11217, 25'd8850, 25'd823, -25'd12452, 25'd6792, -25'd9468, -25'd3808}, '{25'd7924, 25'd2573, -25'd11115, 25'd9159, -25'd9056, 25'd10600, 25'd9880, -25'd3190, -25'd10806}, '{-25'd2779, 25'd11012, -25'd8645, 25'd6278, -25'd8130, 25'd8645, 25'd5763, -25'd4528, -25'd9262}}},
    '{'{'{-25'd1466, 25'd6880, -25'd1128, 25'd11166, 25'd226, 25'd5527, 25'd2256, 25'd1917, -25'd10151}, '{-25'd902, -25'd1128, -25'd8798, 25'd1015, -25'd1015, -25'd4173, -25'd7219, 25'd9926, 25'd7331}, '{-25'd4850, -25'd5752, 25'd4963, 25'd9587, 25'd5188, 25'd10151, -25'd226, 25'd9249, -25'd7219}, '{-25'd7219, 25'd9023, -25'd9813, -25'd2933, -25'd4512, 25'd9700, -25'd1354, 25'd3384, -25'd9926}, '{25'd2707, 25'd1917, -25'd9475, 25'd6655, 25'd5752, -25'd7444, -25'd5414, 25'd3045, -25'd11054}, '{25'd5301, 25'd2030, 25'd7219, 25'd10264, -25'd338, 25'd8121, -25'd2030, 25'd1579, -25'd2143}, '{25'd11392, -25'd8008, -25'd2707, 25'd8911, 25'd2143, -25'd12069, -25'd11843, 25'd9249, -25'd4737}, '{-25'd1354, 25'd4286, -25'd11505, 25'd1692, 25'd1917, 25'd3722, -25'd5188, -25'd2481, 25'd2820}, '{25'd7783, -25'd4061, 25'd3158, -25'd5301, -25'd9136, 25'd6429, -25'd1917, 25'd6316, -25'd902}}, '{'{-25'd9023, 25'd2256, 25'd6993, -25'd8911, -25'd5752, 25'd9023, -25'd5076, -25'd10264, 25'd3497}, '{-25'd11956, -25'd6316, 25'd10151, -25'd8347, -25'd4624, 25'd5978, 25'd9475, -25'd1128, -25'd9587}, '{25'd6542, 25'd9587, 25'd3835, -25'd1015, 25'd9249, 25'd2820, 25'd3722, 25'd10151, 25'd7331}, '{25'd6091, 25'd7783, 25'd6091, -25'd1692, -25'd8459, -25'd4061, -25'd1128, 25'd6316, -25'd2481}, '{25'd11166, -25'd3045, -25'd8121, -25'd9926, -25'd5188, -25'd8347, -25'd11505, -25'd113, -25'd8347}, '{-25'd5076, -25'd8121, 25'd9362, 25'd7444, 25'd4061, -25'd4512, 25'd3835, 25'd1354, -25'd8347}, '{-25'd7106, 25'd0, 25'd7783, 25'd2030, -25'd10151, 25'd6993, 25'd4173, -25'd3158, 25'd2030}, '{25'd4061, 25'd3835, 25'd3497, -25'd1241, -25'd2707, -25'd677, -25'd9813, -25'd1579, -25'd10490}, '{25'd3158, -25'd11730, 25'd677, 25'd4286, 25'd5188, 25'd8008, -25'd8572, -25'd4399, 25'd8347}}, '{'{25'd7331, 25'd10490, -25'd2481, -25'd3497, -25'd5076, 25'd10715, 25'd10602, -25'd2143, 25'd3271}, '{25'd11279, 25'd8008, -25'd677, -25'd2594, -25'd5978, -25'd5978, 25'd1805, -25'd5978, -25'd6429}, '{-25'd1692, 25'd7219, -25'd4399, 25'd12971, 25'd14325, 25'd3045, -25'd6429, 25'd8572, 25'd2594}, '{-25'd3271, 25'd3045, -25'd9136, 25'd2820, -25'd3835, -25'd5188, 25'd12520, 25'd677, -25'd226}, '{25'd6880, 25'd3497, -25'd3271, -25'd4286, 25'd2707, -25'd10038, -25'd6993, -25'd6993, 25'd2707}, '{25'd11279, 25'd3384, 25'd11505, 25'd677, 25'd564, -25'd3948, -25'd10151, 25'd5978, -25'd5414}, '{-25'd7444, 25'd10151, 25'd4737, 25'd3835, -25'd1354, 25'd1015, -25'd677, -25'd10602, -25'd3045}, '{-25'd902, -25'd4737, -25'd451, 25'd7444, -25'd8685, 25'd9475, 25'd5752, 25'd10941, 25'd3384}, '{25'd5865, -25'd8798, 25'd1015, 25'd8459, 25'd8347, 25'd10377, -25'd9362, -25'd11505, 25'd1241}}},
    '{'{'{25'd969, 25'd2787, 25'd4969, -25'd1091, 25'd2787, 25'd9210, 25'd11755, 25'd6665, 25'd1697}, '{25'd7029, 25'd8362, 25'd2424, 25'd14421, 25'd6302, 25'd10422, -25'd4969, -25'd4363, -25'd6786}, '{-25'd6302, 25'd1212, 25'd727, 25'd6059, 25'd7998, -25'd8847, 25'd8968, 25'd2545, -25'd2060}, '{25'd9331, 25'd969, 25'd1575, 25'd6786, 25'd12846, -25'd3151, -25'd7029, 25'd9210, -25'd4847}, '{-25'd5211, 25'd11391, -25'd1697, -25'd6786, -25'd3393, -25'd3757, 25'd2787, 25'd9574, -25'd1939}, '{25'd9574, 25'd727, -25'd7029, -25'd9695, -25'd5938, -25'd5575, -25'd10543, 25'd3030, -25'd12361}, '{25'd9695, 25'd3636, -25'd9816, -25'd7029, -25'd10907, -25'd14785, -25'd3514, -25'd969, -25'd6059}, '{-25'd5332, -25'd9937, 25'd6786, -25'd9695, -25'd13452, 25'd3393, -25'd15512, 25'd4969, -25'd11270}, '{25'd11270, -25'd4241, 25'd8847, 25'd8483, -25'd10058, -25'd1091, -25'd4120, 25'd9937, -25'd4605}}, '{'{25'd1575, 25'd242, 25'd7756, -25'd848, -25'd2666, -25'd8362, -25'd3636, 25'd8483, 25'd485}, '{25'd7998, 25'd9937, -25'd5696, 25'd2545, -25'd1818, 25'd2303, -25'd7998, 25'd4726, -25'd1212}, '{25'd2545, 25'd9574, -25'd2545, -25'd11876, 25'd6665, 25'd8119, 25'd9331, 25'd1091, 25'd3636}, '{25'd4363, 25'd10058, 25'd5332, 25'd606, -25'd8968, -25'd11634, 25'd4605, -25'd7029, -25'd11513}, '{25'd606, 25'd8604, 25'd8968, 25'd8483, -25'd3878, 25'd7877, 25'd7877, -25'd7756, 25'd1091}, '{-25'd11876, -25'd2666, 25'd2424, 25'd4484, 25'd6302, -25'd3393, -25'd8483, 25'd5696, -25'd1575}, '{-25'd2424, 25'd5211, 25'd5938, 25'd1212, 25'd4726, -25'd15148, -25'd3514, 25'd1575, -25'd11634}, '{-25'd8725, 25'd364, -25'd14542, 25'd3272, -25'd7877, 25'd7150, -25'd5696, -25'd5817, 25'd1333}, '{-25'd5938, 25'd9452, 25'd5696, 25'd6544, 25'd364, 25'd5211, 25'd6544, -25'd1212, -25'd11513}}, '{'{-25'd2666, 25'd12240, -25'd3514, -25'd2181, 25'd10422, -25'd10058, 25'd4605, 25'd7271, 25'd6908}, '{25'd2424, 25'd12240, 25'd12724, 25'd3999, -25'd4363, -25'd7877, -25'd4847, 25'd11270, -25'd5817}, '{-25'd242, 25'd3757, 25'd2181, 25'd10907, 25'd9695, 25'd6059, 25'd848, -25'd7029, -25'd3514}, '{-25'd5575, 25'd14663, -25'd3636, 25'd10907, -25'd6665, 25'd7271, -25'd2666, -25'd3272, 25'd10543}, '{25'd4363, 25'd727, 25'd1212, -25'd3272, -25'd7998, -25'd4726, 25'd8241, -25'd10422, 25'd6544}, '{-25'd6302, 25'd12119, -25'd2060, 25'd12603, -25'd7998, 25'd2181, -25'd10785, 25'd4847, -25'd3636}, '{-25'd7756, -25'd8725, 25'd9937, -25'd3030, 25'd10058, -25'd8725, -25'd9210, -25'd3878, -25'd3514}, '{25'd8119, -25'd4484, 25'd7392, 25'd7635, -25'd4969, 25'd9695, -25'd5332, -25'd6059, 25'd8483}, '{-25'd7635, -25'd7513, 25'd9452, -25'd5090, 25'd11391, -25'd3757, -25'd12361, -25'd4484, -25'd13088}}},
    '{'{'{25'd2385, -25'd12469, -25'd9325, -25'd8349, 25'd2060, -25'd6397, 25'd1193, -25'd3578, 25'd10626}, '{25'd6289, 25'd6506, 25'd2385, 25'd2494, 25'd1626, 25'd10409, 25'd0, -25'd9325, -25'd7048}, '{-25'd11494, -25'd11168, -25'd108, 25'd6181, -25'd6397, 25'd4663, 25'd5422, 25'd759, -25'd10518}, '{-25'd10843, 25'd6289, 25'd7915, -25'd6289, 25'd5530, -25'd4771, -25'd7590, 25'd5313, -25'd9542}, '{25'd4554, -25'd10409, -25'd542, 25'd11602, -25'd2385, -25'd3470, -25'd8024, 25'd1843, 25'd7915}, '{-25'd9976, 25'd5855, 25'd9542, 25'd10843, -25'd10951, 25'd5096, -25'd8783, -25'd542, -25'd8458}, '{25'd0, 25'd4879, 25'd10301, -25'd9217, -25'd1735, 25'd1952, 25'd9108, 25'd4771, 25'd12578}, '{25'd11060, -25'd5964, 25'd8891, -25'd3578, 25'd12469, -25'd3036, 25'd217, 25'd12361, 25'd5096}, '{25'd2711, 25'd1735, -25'd10518, 25'd4120, -25'd2277, -25'd3036, -25'd6072, 25'd12253, -25'd4229}}, '{'{-25'd9542, 25'd13337, 25'd11602, 25'd9000, 25'd6723, -25'd2819, -25'd2060, 25'd13228, -25'd4663}, '{25'd5638, -25'd4337, -25'd2928, 25'd7373, 25'd10518, -25'd1735, -25'd3903, 25'd5313, 25'd4879}, '{25'd3253, 25'd651, 25'd10518, 25'd11819, 25'd8241, -25'd867, 25'd976, -25'd9650, 25'd4988}, '{-25'd6614, -25'd8132, 25'd8024, 25'd5205, -25'd542, 25'd9542, -25'd325, 25'd12253, 25'd12578}, '{-25'd5530, 25'd5205, 25'd9000, 25'd3687, 25'd4879, -25'd1193, 25'd7590, 25'd12361, -25'd2602}, '{25'd6723, -25'd8891, 25'd7156, 25'd12686, -25'd3470, 25'd11819, 25'd10192, -25'd8349, 25'd8783}, '{25'd13771, 25'd6614, -25'd5530, 25'd4012, 25'd5096, 25'd9650, -25'd5205, -25'd8674, 25'd8891}, '{25'd7156, 25'd1843, 25'd4988, 25'd7373, -25'd4337, 25'd4012, 25'd3361, 25'd542, 25'd9650}, '{-25'd4771, -25'd3361, 25'd12361, 25'd3578, 25'd10735, -25'd10518, 25'd5313, 25'd2928, -25'd4337}}, '{'{-25'd8566, 25'd6506, -25'd3470, 25'd6397, -25'd9650, -25'd6181, 25'd11060, 25'd1843, 25'd7156}, '{-25'd5313, 25'd12253, 25'd3253, 25'd1735, 25'd3470, -25'd8241, -25'd8458, 25'd1626, 25'd3361}, '{-25'd2819, 25'd2385, 25'd2169, -25'd3036, -25'd1193, -25'd7699, -25'd5747, -25'd4771, 25'd9542}, '{-25'd7265, 25'd3795, 25'd4771, -25'd1193, -25'd1735, -25'd6289, -25'd5530, 25'd6831, -25'd5096}, '{-25'd1843, 25'd10192, 25'd2819, -25'd1301, -25'd434, -25'd4337, -25'd4120, -25'd8349, 25'd7807}, '{25'd2169, -25'd6181, 25'd7048, -25'd4337, -25'd7699, 25'd2928, -25'd1843, -25'd7590, -25'd9325}, '{-25'd5422, -25'd4446, -25'd1626, 25'd8024, -25'd10084, -25'd7807, 25'd7590, -25'd10301, -25'd11385}, '{25'd9325, -25'd6181, -25'd8349, 25'd3903, 25'd976, 25'd3361, 25'd11710, 25'd5747, 25'd6397}, '{-25'd9542, -25'd1843, -25'd9759, -25'd7048, -25'd9325, -25'd2602, 25'd6289, 25'd3795, 25'd3361}}},
    '{'{'{-25'd2359, 25'd1930, -25'd322, -25'd4717, -25'd9220, -25'd4396, -25'd7826, 25'd12972, 25'd9756}, '{25'd7397, -25'd5039, 25'd4074, -25'd6969, 25'd4717, -25'd2680, -25'd536, -25'd8362, -25'd3752}, '{-25'd6111, 25'd7826, 25'd10721, 25'd5039, -25'd4288, 25'd9649, 25'd9970, -25'd214, -25'd4396}, '{-25'd10185, -25'd9434, -25'd3752, 25'd643, 25'd643, -25'd5039, -25'd7719, -25'd4717, -25'd5897}, '{-25'd2787, -25'd2466, 25'd1179, -25'd1930, 25'd9542, 25'd8148, 25'd6969, 25'd5253, -25'd1501}, '{25'd1930, 25'd8362, 25'd7183, -25'd6754, 25'd6969, 25'd3216, -25'd9113, 25'd9327, -25'd4181}, '{25'd7076, 25'd0, 25'd9434, -25'd9113, 25'd6540, 25'd1501, 25'd10399, 25'd214, 25'd7076}, '{-25'd1179, 25'd3323, -25'd3216, -25'd322, -25'd6969, 25'd1823, 25'd1287, 25'd11364, 25'd9970}, '{-25'd536, 25'd5897, 25'd5789, 25'd8470, 25'd3538, -25'd9542, -25'd7719, 25'd9756, 25'd11364}}, '{'{-25'd9542, -25'd11043, -25'd6111, 25'd965, -25'd5897, -25'd965, 25'd1715, -25'd3645, 25'd3860}, '{25'd858, 25'd7933, -25'd13294, 25'd1608, -25'd965, -25'd9327, 25'd6647, -25'd7933, 25'd5146}, '{-25'd6004, 25'd1072, 25'd3109, -25'd1930, -25'd1394, -25'd1823, -25'd8362, 25'd11150, -25'd7076}, '{25'd2251, 25'd4717, 25'd9113, 25'd9327, 25'd4288, -25'd8148, 25'd214, -25'd10292, -25'd9649}, '{-25'd3752, -25'd2037, 25'd1072, 25'd10614, -25'd11579, -25'd7826, -25'd5897, -25'd9113, -25'd5146}, '{25'd1501, 25'd4610, 25'd10935, -25'd6969, -25'd8041, -25'd2466, 25'd2680, -25'd643, 25'd6325}, '{25'd1715, -25'd7933, 25'd4610, 25'd5360, 25'd5789, -25'd536, -25'd6647, -25'd965, -25'd7183}, '{-25'd4610, -25'd9756, -25'd3323, 25'd8148, 25'd214, 25'd3002, 25'd1608, -25'd3109, 25'd1608}, '{25'd7826, 25'd6540, -25'd322, -25'd11257, 25'd7612, 25'd11793, 25'd5575, -25'd858, 25'd2680}}, '{'{-25'd1394, 25'd536, -25'd3216, 25'd1715, -25'd4717, -25'd9113, -25'd6540, 25'd5146, 25'd7933}, '{25'd2466, 25'd6433, -25'd429, -25'd6433, 25'd3752, -25'd8470, 25'd3002, -25'd10399, 25'd4288}, '{-25'd6433, -25'd7505, -25'd2251, -25'd12436, 25'd107, 25'd2895, -25'd11150, 25'd8577, -25'd5146}, '{25'd9542, -25'd965, -25'd7826, -25'd7076, -25'd7612, -25'd1930, -25'd4717, -25'd8041, 25'd5253}, '{-25'd6969, 25'd1287, 25'd5360, -25'd11364, 25'd214, -25'd9649, 25'd0, -25'd5360, -25'd1072}, '{25'd13294, 25'd6969, -25'd5789, 25'd965, 25'd8791, 25'd4503, 25'd6754, -25'd6111, 25'd11471}, '{25'd4288, -25'd4181, -25'd2680, 25'd12543, 25'd5897, -25'd9434, -25'd6540, 25'd13616, 25'd2680}, '{25'd9970, -25'd4610, 25'd6004, -25'd1930, -25'd5253, 25'd12543, -25'd2466, 25'd9756, 25'd6111}, '{25'd8255, 25'd4610, -25'd3323, -25'd1823, 25'd7290, -25'd7933, 25'd7183, 25'd11686, -25'd750}}},
    '{'{'{-25'd5765, 25'd10723, -25'd3690, 25'd7956, -25'd1499, -25'd9109, 25'd115, -25'd6803, -25'd11069}, '{-25'd10377, 25'd1038, -25'd346, 25'd4958, 25'd0, 25'd6342, -25'd1730, -25'd3690, 25'd5304}, '{-25'd4958, 25'd2537, -25'd9455, 25'd2421, -25'd11992, 25'd5535, 25'd1960, -25'd4727, -25'd10839}, '{25'd11069, -25'd1960, -25'd6226, 25'd10147, 25'd8532, -25'd3344, 25'd8994, 25'd4843, 25'd7841}, '{-25'd1614, -25'd2537, 25'd9916, 25'd9570, -25'd8532, 25'd5765, 25'd11069, 25'd5650, -25'd3113}, '{-25'd2421, -25'd9455, -25'd2767, 25'd7149, 25'd1499, 25'd9686, 25'd115, 25'd6457, -25'd8302}, '{25'd7264, 25'd0, -25'd11415, 25'd5765, -25'd2191, 25'd3344, -25'd8071, 25'd8071, 25'd8648}, '{25'd7610, 25'd922, -25'd7264, 25'd3574, -25'd10608, -25'd2075, 25'd346, 25'd10954, -25'd7034}, '{25'd7379, 25'd4497, -25'd1384, 25'd4727, -25'd6457, 25'd10723, -25'd11300, -25'd8417, 25'd6572}}, '{'{25'd7610, -25'd4497, 25'd5419, 25'd9686, -25'd7495, 25'd8302, 25'd4958, 25'd5535, -25'd7610}, '{-25'd3344, -25'd4727, -25'd7034, 25'd346, -25'd7495, -25'd9340, -25'd4958, -25'd9801, -25'd7956}, '{25'd11069, -25'd9109, -25'd692, -25'd4958, -25'd3113, -25'd9686, 25'd11761, 25'd0, 25'd9801}, '{25'd8071, -25'd10262, -25'd577, 25'd10377, -25'd7034, -25'd10954, 25'd7495, 25'd7264, -25'd11184}, '{-25'd461, -25'd3574, 25'd3459, -25'd6457, 25'd4151, 25'd2652, 25'd12107, 25'd2537, -25'd8763}, '{-25'd8763, 25'd5535, -25'd4843, -25'd4151, -25'd5073, 25'd11415, 25'd11761, 25'd1153, -25'd10262}, '{25'd7841, -25'd1153, 25'd11184, 25'd10493, 25'd11069, 25'd9686, 25'd10954, -25'd4382, 25'd1614}, '{25'd6457, 25'd1499, 25'd7841, -25'd692, 25'd9455, -25'd8763, -25'd3229, 25'd1614, -25'd1614}, '{25'd692, -25'd7725, -25'd3229, 25'd6457, -25'd2883, 25'd9916, 25'd7034, -25'd4958, -25'd4266}}, '{'{-25'd6688, -25'd5765, -25'd3574, 25'd1960, -25'd922, -25'd8878, 25'd3690, -25'd2652, -25'd7379}, '{-25'd6918, -25'd6688, 25'd8302, 25'd7956, -25'd12453, -25'd692, 25'd346, -25'd1038, -25'd346}, '{-25'd3113, -25'd4958, -25'd9340, 25'd2767, 25'd6918, 25'd7264, -25'd6226, -25'd2998, 25'd2191}, '{-25'd2421, 25'd231, -25'd12222, 25'd9916, 25'd6572, 25'd8878, -25'd1845, -25'd8532, 25'd7379}, '{25'd5650, -25'd2998, -25'd11876, -25'd3113, -25'd5881, 25'd1038, -25'd8071, 25'd577, -25'd2421}, '{-25'd11300, 25'd4843, 25'd10377, 25'd5996, 25'd6688, -25'd5881, 25'd9916, 25'd10031, 25'd7956}, '{25'd6572, 25'd4382, -25'd3344, 25'd10262, -25'd1499, 25'd4727, 25'd10839, 25'd10608, 25'd9340}, '{-25'd7379, 25'd2883, -25'd7149, -25'd2652, 25'd231, 25'd6342, 25'd10377, -25'd461, 25'd8071}, '{-25'd5650, -25'd10493, 25'd6457, -25'd807, -25'd1153, -25'd8417, -25'd1153, 25'd8648, -25'd14759}}},
    '{'{'{-25'd10363, -25'd8528, 25'd7124, 25'd5613, -25'd11442, -25'd7340, 25'd7988, -25'd9715, -25'd8204}, '{-25'd7232, 25'd2915, -25'd4102, 25'd432, -25'd6908, 25'd8528, 25'd2267, -25'd11658, 25'd3130}, '{25'd4858, 25'd432, 25'd9067, -25'd7232, -25'd12090, 25'd1511, -25'd1619, 25'd9931, 25'd1943}, '{-25'd8851, -25'd5073, 25'd5397, 25'd4750, -25'd3670, 25'd972, 25'd9607, -25'd4750, -25'd10039}, '{25'd2051, -25'd1511, -25'd8204, 25'd3886, 25'd2915, 25'd11010, -25'd216, 25'd2591, -25'd4965}, '{25'd4210, -25'd8096, -25'd7232, -25'd11118, -25'd2267, 25'd1835, -25'd7988, -25'd10902, -25'd10579}, '{-25'd7124, -25'd7988, 25'd2483, -25'd4858, 25'd4210, 25'd972, -25'd5289, -25'd2699, -25'd8204}, '{-25'd5397, -25'd9607, 25'd5289, 25'd7232, -25'd7124, -25'd8096, -25'd7448, -25'd324, -25'd10471}, '{25'd1187, -25'd4210, -25'd4210, 25'd9067, 25'd3238, 25'd1295, -25'd12306, 25'd8312, 25'd5613}}, '{'{25'd6801, -25'd6045, 25'd11010, 25'd1619, -25'd6693, 25'd9715, 25'd12738, -25'd2807, -25'd648}, '{25'd1619, 25'd11658, 25'd7880, 25'd1403, 25'd2699, -25'd2591, 25'd7016, -25'd8096, 25'd3238}, '{-25'd3130, 25'd10687, -25'd7340, -25'd7232, 25'd11442, 25'd4750, 25'd6261, -25'd8636, 25'd7232}, '{25'd0, 25'd7664, -25'd7664, 25'd3022, 25'd6801, -25'd5181, 25'd5721, 25'd7124, -25'd5289}, '{-25'd4965, 25'd7880, 25'd7664, -25'd540, 25'd4965, 25'd11334, -25'd9931, 25'd3562, 25'd5289}, '{25'd13169, 25'd7340, 25'd9283, 25'd108, -25'd4642, 25'd3454, -25'd7664, -25'd2807, 25'd9715}, '{-25'd8312, -25'd972, 25'd2591, -25'd216, -25'd6477, -25'd2375, -25'd10902, -25'd5289, 25'd4102}, '{-25'd3778, -25'd8420, 25'd216, 25'd10579, -25'd1511, 25'd7988, -25'd10039, 25'd10471, 25'd10795}, '{-25'd4102, -25'd9823, 25'd4318, 25'd11874, 25'd7016, 25'd10039, -25'd2591, 25'd10255, 25'd8744}}, '{'{25'd8204, 25'd2807, -25'd108, -25'd8744, -25'd3562, 25'd6908, -25'd1511, -25'd8312, -25'd5829}, '{25'd3454, -25'd7232, 25'd13061, 25'd6369, -25'd2483, 25'd2051, -25'd3562, 25'd9067, 25'd8096}, '{25'd9499, -25'd6045, -25'd1187, 25'd8744, 25'd3454, -25'd9715, -25'd8851, -25'd7664, -25'd3022}, '{25'd10795, 25'd5181, 25'd3994, -25'd3562, 25'd9823, -25'd2591, -25'd9823, 25'd7448, 25'd4858}, '{25'd5613, 25'd2483, -25'd3022, -25'd7340, 25'd3562, 25'd4965, 25'd7556, -25'd5289, 25'd5829}, '{25'd9391, 25'd3886, 25'd5613, 25'd4858, 25'd7664, 25'd1295, -25'd5181, -25'd1943, 25'd6153}, '{-25'd7772, 25'd13709, 25'd5829, 25'd12845, -25'd6045, -25'd6477, -25'd2051, 25'd3022, 25'd1079}, '{25'd7016, -25'd4426, 25'd12630, 25'd1295, -25'd432, 25'd3238, -25'd2267, -25'd6585, 25'd756}, '{25'd10687, 25'd11658, 25'd756, -25'd6477, 25'd3346, -25'd7448, 25'd8420, 25'd12306, -25'd3346}}},
    '{'{'{-25'd3114, 25'd1713, 25'd13548, 25'd6385, -25'd934, -25'd3270, 25'd3114, -25'd4983, 25'd6229}, '{-25'd18842, -25'd3582, 25'd11056, 25'd9188, 25'd11679, 25'd779, -25'd3114, 25'd10745, -25'd9032}, '{-25'd934, -25'd16351, -25'd8565, -25'd12925, -25'd5450, -25'd6385, 25'd9966, 25'd9811, 25'd2803}, '{-25'd8409, 25'd4672, 25'd11368, 25'd7942, -25'd4360, -25'd5295, 25'd13081, -25'd7163, -25'd3270}, '{-25'd2959, 25'd8098, -25'd6073, -25'd8253, 25'd5450, 25'd11523, 25'd7163, 25'd2492, -25'd4672}, '{-25'd9188, -25'd9811, -25'd10589, -25'd3426, -25'd9188, 25'd11991, -25'd8253, -25'd8098, 25'd3582}, '{-25'd7475, 25'd10589, -25'd2647, -25'd1557, -25'd1246, 25'd11991, -25'd5917, -25'd4672, 25'd3426}, '{-25'd5762, -25'd5762, 25'd8876, -25'd1090, 25'd2492, -25'd9188, 25'd2803, -25'd5606, -25'd4516}, '{25'd18220, 25'd4983, 25'd10901, -25'd6540, 25'd12302, -25'd467, -25'd4672, -25'd10901, -25'd11835}}, '{'{-25'd18842, -25'd5762, 25'd7786, -25'd3426, -25'd7475, -25'd11991, 25'd10433, 25'd4516, -25'd11835}, '{-25'd18220, -25'd19933, -25'd8098, 25'd1402, -25'd8876, -25'd12458, -25'd6229, -25'd6696, -25'd9499}, '{-25'd19933, -25'd19933, -25'd11991, -25'd11835, -25'd17752, -25'd3893, 25'd2336, 25'd5139, 25'd5762}, '{25'd5295, 25'd8253, -25'd9811, -25'd7163, -25'd5295, 25'd311, 25'd9188, -25'd3737, -25'd10122}, '{-25'd467, -25'd7942, 25'd12614, 25'd7630, -25'd3582, -25'd2180, -25'd1713, 25'd9966, 25'd3270}, '{-25'd12146, -25'd2492, 25'd1090, 25'd3737, 25'd13236, 25'd10745, 25'd2803, 25'd0, 25'd1713}, '{25'd4827, -25'd3893, 25'd1713, -25'd2336, -25'd3737, 25'd11368, 25'd2180, -25'd9188, 25'd2336}, '{-25'd10122, 25'd6540, 25'd4672, 25'd6540, 25'd10122, -25'd311, 25'd1557, -25'd2336, -25'd1869}, '{25'd5295, 25'd9655, -25'd3270, -25'd8876, -25'd8565, 25'd3737, -25'd3737, -25'd9343, -25'd4049}}, '{'{-25'd18687, -25'd12458, -25'd10745, -25'd3737, 25'd6540, -25'd11679, 25'd2492, 25'd6385, -25'd14482}, '{-25'd12925, -25'd1869, -25'd18220, -25'd5606, -25'd8565, 25'd7008, -25'd9655, 25'd2336, 25'd3426}, '{-25'd19933, -25'd13236, -25'd7786, -25'd14482, 25'd6696, 25'd6696, -25'd1869, -25'd14949, -25'd6073}, '{-25'd3270, -25'd7319, -25'd6229, -25'd10745, -25'd11368, -25'd12458, 25'd5606, -25'd3114, -25'd8409}, '{25'd5450, 25'd1402, 25'd5606, -25'd4049, 25'd7008, -25'd10278, -25'd6229, -25'd11212, -25'd4827}, '{-25'd7942, 25'd6540, -25'd11056, -25'd11056, -25'd3737, -25'd11991, -25'd11991, 25'd7786, -25'd3737}, '{-25'd7942, 25'd934, 25'd5606, 25'd5917, 25'd7319, 25'd5295, -25'd4049, 25'd2959, 25'd6229}, '{25'd3114, 25'd7319, -25'd4049, -25'd11368, -25'd12769, 25'd2180, -25'd6852, 25'd5450, -25'd1869}, '{25'd15417, -25'd1869, -25'd7942, 25'd7008, 25'd7786, -25'd8098, 25'd6229, -25'd13081, 25'd3893}}},
    '{'{'{25'd5726, -25'd487, 25'd12305, 25'd13523, 25'd1827, 25'd5604, -25'd9137, 25'd5117, 25'd7188}, '{25'd2558, 25'd9381, -25'd4630, 25'd5604, 25'd9016, -25'd5970, -25'd8772, -25'd2071, -25'd5239}, '{25'd731, 25'd3046, -25'd2802, -25'd5482, 25'd6944, 25'd5726, -25'd365, -25'd2558, -25'd5482}, '{-25'd6823, 25'd14133, 25'd9625, 25'd8528, -25'd4142, -25'd5482, 25'd5726, 25'd3533, -25'd3655}, '{25'd10478, 25'd8041, 25'd2315, 25'd2437, 25'd9747, -25'd3046, -25'd1218, -25'd5482, 25'd5117}, '{25'd12305, 25'd5482, 25'd5482, 25'd1584, -25'd4751, -25'd6823, -25'd9381, -25'd5848, 25'd975}, '{25'd6701, -25'd4995, -25'd1584, 25'd6335, 25'd10478, -25'd5117, -25'd5239, 25'd4751, 25'd365}, '{25'd14011, -25'd4995, -25'd1706, -25'd5848, 25'd2437, 25'd8041, 25'd8894, 25'd6579, -25'd3777}, '{25'd5604, 25'd13767, -25'd10112, 25'd7310, 25'd4508, 25'd4508, 25'd4142, 25'd9381, -25'd13158}}, '{'{25'd5970, -25'd12671, 25'd244, 25'd7919, -25'd11696, -25'd4020, 25'd975, 25'd8772, 25'd9137}, '{-25'd2924, 25'd3899, 25'd8772, 25'd9625, 25'd2193, 25'd853, -25'd3777, 25'd12671, 25'd122}, '{-25'd975, -25'd2193, -25'd4142, -25'd10843, -25'd487, -25'd7432, -25'd3533, 25'd9747, -25'd4386}, '{-25'd12183, -25'd8772, -25'd1096, -25'd6213, -25'd11818, -25'd3655, -25'd1462, 25'd3899, -25'd7188}, '{-25'd1218, -25'd1462, 25'd3046, -25'd7188, 25'd4751, 25'd7675, -25'd3168, 25'd9990, -25'd853}, '{25'd2680, 25'd0, -25'd10478, 25'd5361, -25'd5970, 25'd8894, 25'd11087, -25'd3533, -25'd9868}, '{25'd487, -25'd12914, -25'd10599, -25'd2315, -25'd4020, -25'd7797, 25'd10599, -25'd9747, 25'd6579}, '{-25'd7188, 25'd7675, 25'd6213, -25'd2924, 25'd3411, 25'd365, -25'd2437, -25'd9381, -25'd9503}, '{-25'd9747, 25'd3168, 25'd122, -25'd244, -25'd6335, 25'd8285, -25'd3046, -25'd8894, -25'd1584}}, '{'{-25'd731, -25'd2680, -25'd4873, -25'd3046, -25'd10234, 25'd4995, -25'd7188, 25'd1949, -25'd1706}, '{-25'd12183, -25'd4142, 25'd6092, -25'd5361, -25'd1218, 25'd4630, -25'd365, 25'd12549, 25'd3411}, '{-25'd11087, -25'd7554, -25'd3411, -25'd5848, 25'd7066, 25'd8894, 25'd7554, 25'd7554, -25'd5117}, '{25'd6579, -25'd15473, 25'd731, -25'd2437, -25'd4630, 25'd3046, 25'd9503, -25'd5361, -25'd5239}, '{-25'd12549, -25'd14011, 25'd1462, 25'd731, -25'd6701, -25'd4995, 25'd7066, 25'd12914, 25'd365}, '{25'd5726, -25'd3046, -25'd8163, -25'd3411, 25'd244, 25'd14985, -25'd2924, 25'd1706, 25'd12792}, '{25'd1340, -25'd10356, 25'd9259, -25'd11696, 25'd4020, -25'd2315, -25'd7310, 25'd9259, 25'd9016}, '{-25'd3411, 25'd4264, -25'd10721, -25'd10721, 25'd9259, -25'd609, -25'd5117, 25'd7919, 25'd11818}, '{-25'd7188, -25'd9503, 25'd8894, 25'd3289, 25'd5361, 25'd6701, -25'd4264, 25'd13402, -25'd6823}}},
    '{'{'{25'd8130, -25'd3786, -25'd3898, -25'd2561, -25'd4566, 25'd11693, -25'd10357, 25'd6459, -25'd10802}, '{25'd2561, -25'd5902, -25'd1448, 25'd7239, 25'd1782, 25'd2673, -25'd557, -25'd6014, -25'd7350}, '{25'd1336, 25'd3675, 25'd891, 25'd2673, 25'd0, -25'd6793, 25'd2561, 25'd2450, -25'd9243}, '{25'd3898, -25'd5791, -25'd3341, 25'd2450, -25'd780, 25'd2005, -25'd1114, -25'd7684, -25'd11582}, '{25'd5680, -25'd7239, 25'd4121, 25'd5011, -25'd4677, 25'd8686, 25'd10914, 25'd6793, -25'd3341}, '{-25'd9800, 25'd111, -25'd3007, -25'd10246, 25'd10023, -25'd4677, -25'd12027, 25'd7239, 25'd1670}, '{-25'd668, 25'd8130, 25'd3786, 25'd223, 25'd1448, 25'd1670, -25'd6682, -25'd8575, -25'd7350}, '{25'd10023, -25'd13030, -25'd1114, -25'd9577, 25'd1559, -25'd7684, 25'd9243, -25'd4677, -25'd12250}, '{-25'd2116, -25'd9021, 25'd1893, 25'd1225, 25'd8018, -25'd2116, -25'd4677, -25'd11359, -25'd1336}}, '{'{25'd0, 25'd7239, -25'd8464, 25'd11805, -25'd7127, 25'd2561, 25'd12807, 25'd6793, 25'd4121}, '{-25'd1225, 25'd2116, 25'd2673, -25'd9021, 25'd8352, -25'd111, -25'd1782, -25'd4900, 25'd12807}, '{25'd5568, 25'd3898, -25'd5568, 25'd780, -25'd7127, 25'd6905, 25'd7461, 25'd12362, -25'd3341}, '{-25'd9021, 25'd7684, -25'd2784, 25'd1336, 25'd6793, -25'd3230, -25'd1225, -25'd6014, 25'd7350}, '{25'd8909, 25'd11248, 25'd10468, 25'd4789, 25'd557, -25'd2005, 25'd9689, 25'd13587, -25'd1782}, '{-25'd334, 25'd4566, -25'd2784, 25'd7350, -25'd5123, -25'd111, 25'd9466, 25'd4789, 25'd4789}, '{-25'd5457, 25'd6682, 25'd7573, -25'd8018, -25'd3341, 25'd13809, 25'd4677, 25'd8798, 25'd14143}, '{-25'd111, -25'd111, -25'd9243, 25'd1114, -25'd7907, 25'd1448, -25'd8018, 25'd3007, 25'd3118}, '{25'd2784, -25'd2005, -25'd6905, -25'd7350, -25'd3118, -25'd3675, 25'd12918, -25'd557, -25'd6236}}, '{'{-25'd10468, -25'd668, -25'd7127, 25'd1559, 25'd10580, 25'd3230, -25'd10134, -25'd111, -25'd2227}, '{-25'd2673, -25'd8018, 25'd1114, 25'd1893, -25'd9689, -25'd8241, 25'd6793, 25'd10134, 25'd10134}, '{-25'd4566, 25'd5568, 25'd2005, 25'd10023, -25'd1559, -25'd7127, 25'd11582, -25'd2450, 25'd7461}, '{-25'd3007, 25'd11248, -25'd7573, -25'd5568, 25'd7796, -25'd111, -25'd10691, -25'd2784, -25'd7684}, '{25'd7796, 25'd7907, -25'd4121, -25'd2116, 25'd5123, 25'd445, -25'd7796, -25'd3118, 25'd9911}, '{-25'd9911, -25'd7684, 25'd1114, 25'd9355, -25'd4900, -25'd5234, -25'd5234, -25'd2227, 25'd6459}, '{25'd1114, -25'd1002, 25'd6793, 25'd11916, 25'd9243, 25'd2784, 25'd1336, -25'd8575, -25'd9466}, '{-25'd1114, -25'd6348, -25'd8575, 25'd2116, -25'd8352, -25'd5902, 25'd0, 25'd10914, 25'd10468}, '{25'd3675, 25'd11805, 25'd2561, 25'd6348, 25'd12473, -25'd3341, 25'd6793, 25'd9466, 25'd3007}}},
    '{'{'{25'd3078, 25'd7035, 25'd10442, 25'd11542, 25'd7585, -25'd7914, -25'd8904, 25'd8024, -25'd8684}, '{25'd7365, 25'd9343, -25'd8354, 25'd9783, -25'd9563, 25'd7255, -25'd4287, -25'd220, -25'd330}, '{25'd4287, 25'd1759, -25'd7694, 25'd3188, -25'd2858, 25'd10113, 25'd4946, 25'd1429, 25'd8354}, '{25'd1319, -25'd8904, -25'd2638, -25'd4946, 25'd7914, -25'd1979, -25'd8464, 25'd110, -25'd7145}, '{25'd8464, 25'd3737, 25'd7255, -25'd6925, -25'd2198, -25'd2198, 25'd3408, -25'd8684, 25'd10552}, '{-25'd8024, 25'd8244, -25'd8134, -25'd6265, 25'd6046, -25'd5276, -25'd879, 25'd6705, 25'd1099}, '{-25'd2968, 25'd7804, 25'd5826, -25'd1979, -25'd769, 25'd2638, -25'd10442, 25'd769, 25'd10772}, '{-25'd1649, 25'd3847, 25'd3078, -25'd11652, -25'd110, 25'd4287, 25'd330, 25'd5826, 25'd1099}, '{25'd6265, -25'd5166, -25'd4946, -25'd1319, 25'd5826, 25'd4397, 25'd1099, 25'd5936, -25'd3737}}, '{'{25'd6156, -25'd2528, -25'd8904, 25'd3517, 25'd11981, 25'd1979, -25'd7145, 25'd989, 25'd1429}, '{25'd2088, 25'd12751, 25'd1429, 25'd6156, -25'd7914, 25'd12091, -25'd8904, -25'd5936, 25'd8354}, '{25'd5716, 25'd3408, 25'd769, 25'd2638, -25'd769, 25'd5826, 25'd12091, 25'd2858, -25'd3847}, '{-25'd7914, 25'd3957, -25'd10113, -25'd6485, 25'd5826, 25'd1099, 25'd3078, 25'd4617, 25'd10772}, '{25'd13960, 25'd8024, 25'd1429, 25'd10552, -25'd5716, 25'd11102, -25'd1429, -25'd4837, 25'd4727}, '{-25'd989, 25'd7365, 25'd6925, -25'd2198, 25'd10662, 25'd10003, 25'd7585, 25'd11212, 25'd330}, '{-25'd3078, 25'd12531, 25'd5606, 25'd9563, 25'd3517, 25'd6265, 25'd8354, 25'd0, -25'd7804}, '{-25'd8574, -25'd2418, 25'd11432, -25'd2308, 25'd12091, 25'd0, -25'd8904, -25'd110, -25'd7585}, '{25'd6595, -25'd440, 25'd220, 25'd7255, -25'd4287, 25'd12531, -25'd3188, 25'd3847, 25'd12641}}, '{'{-25'd6485, -25'd1869, -25'd5716, 25'd1649, -25'd10223, 25'd4837, -25'd13630, -25'd13520, -25'd13191}, '{-25'd7585, -25'd2198, -25'd10772, 25'd6705, 25'd7694, 25'd1979, 25'd4727, -25'd7145, 25'd1319}, '{-25'd2638, -25'd7585, 25'd7255, -25'd3737, 25'd8354, -25'd12201, -25'd12641, 25'd8134, -25'd11542}, '{25'd5386, 25'd3737, -25'd5166, -25'd3737, -25'd1979, 25'd5496, 25'd3627, -25'd10662, 25'd989}, '{25'd4727, 25'd2088, 25'd8574, 25'd7475, -25'd11981, -25'd4287, -25'd11981, 25'd8574, -25'd8574}, '{-25'd2088, 25'd6265, -25'd4177, -25'd9673, -25'd9233, -25'd3078, -25'd3847, 25'd7475, -25'd660}, '{-25'd6485, 25'd10003, 25'd11322, -25'd769, -25'd3847, -25'd1209, 25'd5056, -25'd6265, 25'd6705}, '{-25'd1099, -25'd10882, -25'd1539, 25'd1209, -25'd5496, -25'd10442, 25'd6595, 25'd7804, -25'd2528}, '{25'd220, -25'd330, -25'd2638, 25'd3627, -25'd3737, -25'd5056, 25'd6705, -25'd5166, 25'd7585}}},
    '{'{'{25'd6608, -25'd1322, -25'd2247, 25'd8458, -25'd6211, 25'd7797, -25'd3965, 25'd10176, -25'd3832}, '{25'd10308, 25'd16784, 25'd6343, 25'd15991, -25'd2114, 25'd1982, 25'd5022, 25'd11233, 25'd7401}, '{25'd7665, -25'd2775, -25'd4890, 25'd6740, 25'd7004, 25'd7004, 25'd2643, -25'd10572, -25'd7929}, '{25'd13215, 25'd11101, 25'd5815, -25'd3436, -25'd10969, 25'd2511, -25'd9119, -25'd264, -25'd8590}, '{-25'd1850, -25'd661, -25'd5022, 25'd396, -25'd7269, -25'd4493, -25'd13612, 25'd5418, -25'd5286}, '{25'd5154, 25'd529, -25'd9515, -25'd2775, 25'd925, -25'd11762, -25'd5683, -25'd14405, 25'd2907}, '{25'd3965, 25'd10572, 25'd4493, -25'd13083, -25'd3304, 25'd5154, -25'd14405, -25'd6740, 25'd529}, '{25'd8722, 25'd4493, 25'd529, 25'd1057, 25'd1850, -25'd529, -25'd12819, -25'd12687, -25'd5947}, '{25'd2907, 25'd3568, -25'd13083, -25'd1454, -25'd7136, -25'd5154, -25'd1850, -25'd7929, -25'd7797}}, '{'{25'd7533, -25'd3172, 25'd1189, -25'd6872, -25'd3436, 25'd264, 25'd7004, 25'd925, 25'd9383}, '{25'd3040, -25'd1586, -25'd3568, 25'd8722, 25'd5551, 25'd5551, 25'd9912, -25'd7533, -25'd1850}, '{25'd11762, 25'd5683, 25'd6608, 25'd8194, 25'd2511, -25'd7797, -25'd7269, 25'd396, -25'd4361}, '{25'd1189, -25'd1718, -25'd4493, -25'd1718, 25'd5022, 25'd4493, -25'd396, -25'd7401, -25'd4493}, '{25'd8722, 25'd5418, -25'd10176, 25'd1322, -25'd3172, 25'd11101, -25'd5815, -25'd3568, 25'd1586}, '{-25'd1322, -25'd9647, -25'd661, -25'd8854, -25'd10572, -25'd9912, 25'd2247, 25'd5551, 25'd8854}, '{-25'd4890, -25'd3965, -25'd4625, -25'd10837, 25'd5551, -25'd1850, -25'd7136, -25'd3304, -25'd2775}, '{25'd3436, -25'd7929, -25'd6343, -25'd11762, 25'd7533, -25'd9251, 25'd4097, 25'd4361, -25'd11894}, '{25'd10044, 25'd5947, 25'd793, -25'd4097, 25'd8458, -25'd6476, 25'd264, -25'd12555, -25'd9779}}, '{'{-25'd4625, -25'd4361, -25'd1057, 25'd4493, 25'd5815, -25'd2114, -25'd132, 25'd13612, -25'd2775}, '{25'd12819, 25'd2511, 25'd0, 25'd5286, -25'd5551, 25'd14405, -25'd396, -25'd6476, 25'd3700}, '{25'd3965, -25'd7004, 25'd4758, -25'd6211, -25'd6343, -25'd7004, 25'd6608, -25'd5154, -25'd8458}, '{-25'd3172, 25'd661, 25'd3965, 25'd793, -25'd3832, 25'd9383, -25'd1718, 25'd6211, 25'd11233}, '{-25'd2643, -25'd6079, 25'd12158, 25'd132, 25'd13083, 25'd1718, -25'd1057, 25'd10837, 25'd1586}, '{25'd14537, 25'd5551, -25'd4625, -25'd1718, -25'd8194, 25'd6079, 25'd7533, 25'd2511, 25'd12951}, '{25'd396, -25'd6872, 25'd4229, -25'd2643, -25'd8326, -25'd10440, -25'd1982, 25'd6608, 25'd3040}, '{25'd10572, 25'd10572, -25'd2247, 25'd396, -25'd1454, 25'd7269, 25'd5947, -25'd9912, -25'd5418}, '{25'd1189, 25'd7401, 25'd1057, -25'd5154, 25'd8854, 25'd2247, -25'd6608, 25'd0, -25'd10572}}},
    '{'{'{25'd9086, -25'd4073, 25'd2715, 25'd9921, 25'd9817, 25'd9190, -25'd6057, 25'd9086, 25'd6579}, '{-25'd11070, -25'd9817, 25'd2506, 25'd1567, -25'd522, 25'd11383, -25'd1044, -25'd5848, 25'd2715}, '{25'd1462, 25'd4804, -25'd4177, -25'd6788, 25'd10443, -25'd313, -25'd4491, -25'd1567, -25'd9921}, '{-25'd7102, 25'd10966, 25'd11488, 25'd9086, -25'd7728, -25'd10861, -25'd4073, -25'd10130, -25'd313}, '{25'd3133, -25'd7102, -25'd835, 25'd10548, 25'd11906, 25'd104, 25'd11488, -25'd7415, 25'd3342}, '{-25'd5117, 25'd10026, 25'd3655, 25'd5013, 25'd6684, -25'd5639, 25'd627, 25'd3446, -25'd1253}, '{25'd11383, 25'd8773, 25'd6057, -25'd4177, 25'd9712, -25'd4491, 25'd10235, 25'd2715, -25'd7102}, '{25'd9608, 25'd10861, -25'd5848, 25'd3551, 25'd4386, -25'd4282, 25'd8355, -25'd1462, -25'd10339}, '{-25'd8877, 25'd10443, -25'd8355, -25'd3655, 25'd7624, 25'd10966, 25'd7310, 25'd8564, 25'd3342}}, '{'{25'd8355, -25'd2924, -25'd9712, 25'd1462, -25'd9817, -25'd5117, 25'd5326, -25'd5639, -25'd10861}, '{25'd7624, 25'd7624, -25'd9712, 25'd7415, 25'd5535, 25'd8146, -25'd12532, -25'd9712, -25'd8564}, '{25'd8459, -25'd11906, 25'd2715, 25'd8041, 25'd418, 25'd2611, -25'd11906, 25'd209, -25'd5639}, '{-25'd9295, 25'd3655, -25'd418, -25'd3237, -25'd5744, -25'd8981, 25'd10548, 25'd2089, 25'd4700}, '{-25'd9504, -25'd10339, -25'd104, 25'd8355, 25'd3655, -25'd5848, -25'd3029, -25'd12741, 25'd9921}, '{-25'd13054, -25'd9921, 25'd5222, -25'd4073, 25'd5222, -25'd7310, 25'd10966, 25'd4908, 25'd731}, '{25'd6997, -25'd13263, -25'd4386, 25'd3760, -25'd10026, 25'd1567, -25'd9921, -25'd2402, -25'd2715}, '{-25'd3342, -25'd5848, 25'd3029, 25'd6893, 25'd4491, -25'd8459, -25'd9921, 25'd2611, 25'd3760}, '{25'd9295, -25'd4804, -25'd731, 25'd1044, 25'd7206, -25'd10235, -25'd1671, -25'd11383, -25'd6371}}, '{'{25'd522, -25'd5744, -25'd7102, -25'd11383, 25'd4700, 25'd8459, 25'd8877, -25'd11175, -25'd8250}, '{-25'd5222, -25'd12114, -25'd418, -25'd2506, 25'd5848, -25'd6057, -25'd10548, -25'd11279, -25'd2611}, '{-25'd10130, -25'd7728, 25'd9086, 25'd5953, 25'd4282, 25'd4073, -25'd3864, 25'd7519, 25'd8564}, '{25'd2402, 25'd3133, -25'd5639, -25'd6893, 25'd1775, -25'd5013, -25'd3864, 25'd104, 25'd3864}, '{-25'd8877, -25'd9817, -25'd4386, 25'd9086, -25'd5744, -25'd7624, -25'd8146, -25'd1253, -25'd1358}, '{25'd9921, 25'd522, -25'd3133, -25'd2924, 25'd2506, 25'd10548, 25'd209, 25'd5431, 25'd7415}, '{-25'd5222, -25'd10443, 25'd522, 25'd4073, -25'd10757, -25'd7937, -25'd313, 25'd209, -25'd9295}, '{25'd7206, -25'd10339, -25'd10861, 25'd8250, 25'd10861, -25'd2402, -25'd8355, -25'd7519, 25'd1462}, '{25'd1044, 25'd3655, -25'd4700, -25'd11175, -25'd10339, 25'd11488, 25'd9086, -25'd9921, 25'd5535}}},
    '{'{'{-25'd4883, -25'd9875, -25'd2062, -25'd1194, 25'd8356, -25'd3255, 25'd3581, 25'd9441, 25'd3798}, '{25'd4775, 25'd10743, 25'd0, -25'd12696, -25'd6402, -25'd7162, -25'd4449, -25'd1411, 25'd4341}, '{25'd7813, -25'd651, 25'd1845, 25'd2387, -25'd12370, -25'd5317, -25'd3364, 25'd9007, 25'd2062}, '{25'd7704, 25'd5751, -25'd7704, 25'd2279, 25'd7596, -25'd10960, 25'd7596, -25'd11394, -25'd7379}, '{-25'd11068, 25'd7487, -25'd12045, 25'd10417, -25'd10743, 25'd10743, 25'd8138, 25'd4123, 25'd12153}, '{-25'd760, -25'd1736, -25'd6185, -25'd4449, -25'd1845, -25'd10200, 25'd2062, -25'd7813, -25'd109}, '{25'd7270, 25'd1736, 25'd7053, -25'd2713, -25'd7813, 25'd8138, 25'd5751, -25'd7270, -25'd6836}, '{-25'd4341, -25'd6728, -25'd10960, 25'd6294, -25'd6294, 25'd3255, 25'd8464, -25'd10200, -25'd6619}, '{25'd7379, 25'd3581, -25'd109, -25'd3038, 25'd3906, 25'd4775, 25'd5317, -25'd2930, 25'd3255}}, '{'{25'd8030, 25'd12588, 25'd2713, -25'd326, 25'd2604, 25'd3472, -25'd5860, 25'd12479, 25'd7704}, '{-25'd5426, -25'd7270, -25'd7162, 25'd2496, 25'd6619, 25'd4558, -25'd1845, 25'd4232, 25'd2930}, '{25'd6185, -25'd8030, -25'd6294, 25'd6511, -25'd9875, 25'd6402, -25'd5317, -25'd8247, -25'd7162}, '{25'd8464, -25'd8247, -25'd5860, -25'd1194, 25'd6511, 25'd11611, 25'd1302, -25'd2604, 25'd4232}, '{-25'd2496, 25'd1519, -25'd1194, 25'd5534, 25'd2930, 25'd2387, -25'd8898, 25'd5751, 25'd3689}, '{25'd13781, 25'd9658, 25'd5534, -25'd8898, 25'd7596, 25'd2496, 25'd7379, -25'd11068, -25'd2170}, '{25'd868, 25'd1845, 25'd1736, 25'd10200, 25'd9766, 25'd5643, -25'd3364, 25'd1411, -25'd5643}, '{-25'd6836, -25'd7379, -25'd5100, 25'd1519, 25'd11068, 25'd4992, -25'd4992, 25'd11068, 25'd6402}, '{25'd3906, -25'd9658, 25'd5426, 25'd2821, 25'd8356, -25'd7704, 25'd3906, -25'd3147, -25'd5860}}, '{'{-25'd9007, 25'd7921, -25'd9007, 25'd8681, 25'd868, -25'd4558, -25'd8464, 25'd4558, 25'd651}, '{-25'd10092, -25'd3798, 25'd6185, 25'd8681, 25'd4666, 25'd9766, 25'd7053, 25'd6619, 25'd8790}, '{-25'd7053, -25'd8138, 25'd9766, 25'd3364, 25'd2604, 25'd8356, -25'd11068, -25'd1953, -25'd4123}, '{25'd1519, -25'd5209, -25'd8247, 25'd6077, 25'd8030, 25'd6619, 25'd5860, 25'd1194, 25'd3906}, '{25'd11719, -25'd434, 25'd0, -25'd8898, -25'd8681, -25'd11285, -25'd4558, 25'd977, 25'd9658}, '{-25'd6077, -25'd10851, 25'd6185, 25'd3147, 25'd8030, -25'd12153, 25'd2387, 25'd543, 25'd4775}, '{-25'd7596, -25'd8573, 25'd9224, 25'd5209, -25'd1736, -25'd11611, 25'd2496, -25'd11285, -25'd4232}, '{25'd6511, 25'd2930, 25'd7813, -25'd7704, 25'd8898, -25'd4123, -25'd1411, -25'd10634, -25'd1519}, '{-25'd217, -25'd5100, -25'd5643, 25'd10200, 25'd8790, 25'd9549, 25'd543, 25'd5534, -25'd4449}}}
};
