localparam bit signed [0:2][0:7][0:2][0:2][19:0] Weight3 = '{
    '{'{'{-20'd524288, 20'd524287, -20'd524288}, '{20'd116063, 20'd464250, 20'd0}, '{-20'd333680, 20'd210363, 20'd65285}}, '{'{-20'd87047, 20'd79793, -20'd311918}, '{-20'd377203, -20'd427981, 20'd43523}, '{20'd87047, 20'd130570, -20'd326426}}, '{'{-20'd72539, 20'd377203, 20'd282902}, '{20'd515027, 20'd224871, 20'd524287}, '{20'd435234, 20'd181348, 20'd174094}}, '{'{20'd515027, -20'd290156, -20'd369949}, '{-20'd524288, -20'd290156, -20'd108809}, '{-20'd166840, -20'd43523, -20'd188602}}, '{'{20'd398965, 20'd435234, 20'd87047}, '{20'd340934, 20'd7254, 20'd188602}, '{20'd253887, -20'd94301, -20'd123316}}, '{'{20'd195856, 20'd152332, -20'd152332}, '{-20'd87047, -20'd145078, 20'd145078}, '{-20'd203109, -20'd275648, 20'd123316}}, '{'{-20'd203109, -20'd246633, -20'd348188}, '{20'd58031, 20'd29016, -20'd181348}, '{20'd304664, 20'd333680, -20'd7254}}, '{'{-20'd152332, 20'd195856, 20'd348188}, '{20'd524287, 20'd217617, -20'd145078}, '{20'd29016, 20'd464250, -20'd7254}}},
    '{'{'{-20'd524288, 20'd524287, -20'd265295}, '{20'd524287, 20'd435841, 20'd9475}, '{-20'd524288, 20'd28424, -20'd350568}}, '{'{-20'd341093, -20'd360043, 20'd217921}, '{-20'd246345, -20'd255820, 20'd85273}, '{-20'd151597, 20'd113698, 20'd94748}}, '{'{-20'd189496, 20'd303194, -20'd104223}, '{-20'd265295, -20'd104223, 20'd75798}, '{20'd274769, 20'd435841, -20'd331618}}, '{'{20'd524287, 20'd208446, -20'd227395}, '{-20'd123172, -20'd132647, 20'd524287}, '{-20'd28424, -20'd274769, 20'd416891}}, '{'{20'd113698, -20'd9475, 20'd397942}, '{-20'd161072, -20'd123172, 20'd161072}, '{20'd303194, 20'd303194, -20'd28424}}, '{'{-20'd236870, 20'd454791, 20'd524287}, '{20'd227395, 20'd227395, 20'd217921}, '{-20'd255820, 20'd37899, 20'd524287}}, '{'{-20'd132647, -20'd331618, -20'd303194}, '{20'd170546, 20'd284244, 20'd312669}, '{20'd94748, -20'd56849, 20'd9475}}, '{'{-20'd56849, 20'd123172, 20'd524287}, '{20'd37899, -20'd161072, -20'd151597}, '{-20'd104223, 20'd360043, 20'd161072}}},
    '{'{'{-20'd515185, 20'd84303, -20'd524288}, '{-20'd524288, -20'd215441, -20'd412148}, '{-20'd524288, 20'd524287, -20'd524288}}, '{'{-20'd149872, -20'd84303, -20'd524288}, '{-20'd28101, -20'd421515, -20'd468350}, '{-20'd524288, -20'd37468, -20'd430882}}, '{'{20'd458983, 20'd74936, 20'd28101}, '{20'd468350, 20'd524287, 20'd421515}, '{-20'd46835, 20'd496451, -20'd37468}}, '{'{20'd65569, 20'd131138, 20'd65569}, '{20'd524287, 20'd271643, 20'd393414}, '{-20'd421515, 20'd56202, 20'd46835}}, '{'{-20'd177973, -20'd65569, 20'd46835}, '{20'd468350, 20'd393414, 20'd505818}, '{20'd524287, 20'd93670, 20'd187340}}, '{'{-20'd140505, -20'd290377, -20'd271643}, '{-20'd365313, -20'd402781, 20'd18734}, '{-20'd449616, 20'd121771, -20'd290377}}, '{'{-20'd9367, 20'd224808, -20'd327845}, '{-20'd159239, -20'd215441, -20'd159239}, '{20'd187340, -20'd9367, -20'd9367}}, '{'{20'd468350, 20'd65569, 20'd131138}, '{20'd159239, -20'd103037, 20'd412148}, '{-20'd112404, 20'd28101, 20'd402781}}}
};
