localparam bit signed [0:26][19:0] Output3 = '{20'd164, 20'd169, 20'd87, 20'd20, -20'd80, 20'd103, 20'd201, -20'd107, -20'd39, 20'd158, 20'd142, -20'd17, -20'd66, -20'd116, 20'd91, -20'd17, 20'd163, -20'd22, -20'd87, -20'd134, -20'd90, -20'd22, -20'd72, -20'd321, 20'd37, 20'd70, -20'd107};
