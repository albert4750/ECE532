logic signed [7:0] layer3_weight[3][12][4][4] = '{
    '{
        '{'{107, -2, 3, -64}, '{-91, 119, 39, -116}, '{-44, 75, -52, -8}, '{-14, 91, 47, -71}},
        '{'{21, -20, -116, 111}, '{17, 39, 31, -17}, '{29, 55, 65, -91}, '{-128, -105, 13, 8}},
        '{'{84, -75, 82, -48}, '{-115, 8, 6, 27}, '{37, 35, -88, 26}, '{-34, 76, 57, -83}},
        '{'{-48, -70, 23, 126}, '{114, 106, 72, 119}, '{118, 80, 117, -3}, '{-110, 74, 15, 102}},
        '{'{-3, -40, 100, 111}, '{-64, 3, 90, 20}, '{111, 47, 62, -31}, '{-104, 82, -88, 9}},
        '{'{-56, 71, 92, 111}, '{-87, -109, 86, -61}, '{119, 78, -1, -9}, '{-62, 87, 107, -104}},
        '{'{-44, 35, -6, 46}, '{-96, -94, -86, -36}, '{-91, 100, -46, -73}, '{-22, -93, 103, -29}},
        '{'{-63, -35, 20, 101}, '{-29, -82, -30, -37}, '{-66, -66, 113, 123}, '{-50, -22, 30, -37}},
        '{'{-77, -124, 68, 6}, '{105, -87, -125, 39}, '{108, -28, 27, 13}, '{-84, -128, -54, 93}},
        '{'{-50, 0, -128, -32}, '{-12, -117, -99, 5}, '{-59, 57, -98, -110}, '{-22, -112, -9, -47}},
        '{'{75, -119, 9, 90}, '{-52, 64, 103, 28}, '{118, -51, -41, 58}, '{-7, 48, 27, -21}},
        '{'{25, 84, -17, -52}, '{-104, -123, -94, -52}, '{59, -85, 79, -69}, '{-107, 100, 113, 126}}
    },
    '{
        '{'{-20, -116, -16, -30}, '{5, -108, -4, 31}, '{-30, -105, -109, -43}, '{-81, 122, -122, -60}},
        '{'{73, -104, 47, 32}, '{74, 90, 91, -112}, '{98, 22, -3, -100}, '{-100, -15, 78, -27}},
        '{'{-39, 5, -62, 35}, '{75, 51, -51, 99}, '{56, 95, 94, -123}, '{-99, -37, 121, 53}},
        '{'{65, -67, 104, 26}, '{-100, 103, 39, -31}, '{-23, 47, -19, 32}, '{-7, -124, 54, 0}},
        '{'{-117, 51, -29, 68}, '{-102, -113, 113, 92}, '{-22, 16, -12, -58}, '{120, -33, -126, 124}},
        '{'{-111, 114, -63, 32}, '{97, 38, -60, -34}, '{-124, 123, -49, -1}, '{-107, -7, -13, -26}},
        '{'{-118, -112, -126, -82}, '{61, 46, -18, -96}, '{103, 23, 61, 1}, '{-92, -39, -120, -81}},
        '{'{-37, -128, 35, -102}, '{62, -17, 52, 106}, '{22, 31, 1, -35}, '{-125, -125, -30, -12}},
        '{'{36, 42, -18, -108}, '{105, 5, 88, 127}, '{-45, 54, 101, -125}, '{-45, 23, -80, -34}},
        '{'{30, 89, 7, 42}, '{12, -124, 112, 27}, '{76, -17, 74, 124}, '{43, 53, 110, 10}},
        '{'{115, -85, -122, 71}, '{-128, -77, 34, -32}, '{-105, 64, 71, 30}, '{-110, -96, -126, 38}},
        '{'{-116, -64, -2, 124}, '{-56, -125, 13, -2}, '{90, 3, 102, 70}, '{6, 20, -70, -126}}
    },
    '{
        '{'{85, 47, 127, 52}, '{-70, -18, -46, 126}, '{-48, -71, 43, -95}, '{106, -59, 93, -49}},
        '{'{-39, 109, 117, -104}, '{-28, 60, -7, -64}, '{61, -51, -116, 70}, '{-15, -79, 3, 32}},
        '{'{-13, 49, 99, 13}, '{-53, -111, -60, 87}, '{-81, -54, 38, -12}, '{117, -26, 48, -92}},
        '{'{93, -103, -93, 71}, '{64, -64, -120, 67}, '{-122, -27, 124, 7}, '{51, 77, -46, -8}},
        '{'{-111, -125, -2, -120}, '{-81, -85, 61, -125}, '{-84, -53, 117, -79}, '{-78, 10, 43, 79}},
        '{'{91, -26, -66, 99}, '{-46, 125, -66, -11}, '{35, -43, 28, 59}, '{97, -39, 74, -127}},
        '{'{122, 21, 25, 10}, '{-8, 41, -115, 51}, '{-62, 82, 84, 7}, '{-88, -72, -43, -91}},
        '{'{46, 83, 90, 55}, '{6, -128, 8, 124}, '{85, -5, 111, 37}, '{67, 46, 104, 41}},
        '{'{-36, -65, -71, 119}, '{-28, -89, 65, 51}, '{61, -19, 69, 58}, '{-37, -33, 40, -55}},
        '{'{53, -8, -121, -29}, '{47, 69, 41, -100}, '{118, -6, -43, -117}, '{-125, -110, 35, -82}},
        '{'{-23, 17, -17, 27}, '{-74, -17, 73, 19}, '{71, -57, -27, 43}, '{126, 44, -18, 46}},
        '{'{34, 33, -54, -9}, '{-59, 92, -82, 32}, '{83, 39, 30, 95}, '{-17, 47, 1, 32}}
    }
};
