logic signed [7:0] convolve4_weight[4][8][3][3] = '{
    '{
        '{'{-4, -11, -28}, '{-38, -60, -23}, '{-118, -116, -24}},
        '{'{97, 37, 39}, '{32, -6, -95}, '{26, -29, 89}},
        '{'{-78, -40, 82}, '{-108, 94, 28}, '{-56, -110, 25}},
        '{'{24, -89, 106}, '{-5, -100, 24}, '{18, 67, 44}},
        '{'{83, -83, -74}, '{-128, 10, 67}, '{6, 91, -29}},
        '{'{57, 70, 19}, '{34, -78, 114}, '{-26, -108, 43}},
        '{'{-10, 0, 100}, '{-19, -23, 66}, '{97, 12, -113}},
        '{'{-10, -95, 23}, '{12, 5, -90}, '{-127, -118, -122}}
    },
    '{
        '{'{-3, -122, -26}, '{38, -53, -14}, '{-43, -2, -14}},
        '{'{50, -77, -126}, '{-52, 29, -119}, '{-13, 72, 5}},
        '{'{-12, 53, 107}, '{65, -85, -49}, '{-66, -52, -81}},
        '{'{-52, 21, -8}, '{-110, -39, -115}, '{94, -36, 108}},
        '{'{-23, 85, -122}, '{-28, -80, -88}, '{26, 30, 5}},
        '{'{15, 63, 101}, '{-91, -69, -15}, '{-33, -32, 112}},
        '{'{80, -96, -66}, '{10, 12, -35}, '{-64, 29, -38}},
        '{'{103, 22, 19}, '{5, -92, -45}, '{-1, 100, -123}}
    },
    '{
        '{'{-36, 76, 26}, '{113, -45, 12}, '{102, 7, 52}},
        '{'{-48, 29, -128}, '{87, 79, -54}, '{124, 3, -67}},
        '{'{-61, 16, -16}, '{73, -44, -12}, '{101, 127, -72}},
        '{'{-66, 56, -80}, '{17, -11, 57}, '{-119, 108, 62}},
        '{'{-49, 102, 78}, '{33, 4, 16}, '{100, -57, -66}},
        '{'{-105, -37, -18}, '{-121, 125, -106}, '{-30, 30, 118}},
        '{'{-48, 27, -81}, '{111, -14, -117}, '{87, -50, 103}},
        '{'{-98, -38, -94}, '{-74, -47, 35}, '{-57, -19, -69}}
    },
    '{
        '{'{-16, 37, -60}, '{53, -115, -27}, '{-109, -21, -120}},
        '{'{-32, 81, 69}, '{-4, -28, 1}, '{125, 29, 5}},
        '{'{80, 102, 120}, '{40, 22, -98}, '{127, -109, -124}},
        '{'{20, -22, -54}, '{-5, 67, 86}, '{-68, 101, 122}},
        '{'{-35, 41, -88}, '{60, 81, 51}, '{-88, -69, 106}},
        '{'{94, -99, 97}, '{-34, 110, 37}, '{-2, 88, -112}},
        '{'{-29, 39, 29}, '{124, -63, -105}, '{72, 0, -41}},
        '{'{-91, -17, 63}, '{26, 89, -39}, '{6, 88, 119}}
    }
};
