localparam bit signed [0:7][0:7][0:2][0:2][24:0] Weight2 = '{
    '{'{'{-25'd5712, -25'd4200, -25'd4536}, '{-25'd8232, -25'd7392, -25'd14448}, '{25'd6720, -25'd336, -25'd5040}}, '{'{25'd168, -25'd1512, 25'd1512}, '{25'd2016, -25'd336, 25'd1176}, '{25'd1344, 25'd1344, 25'd2856}}, '{'{25'd8064, 25'd6384, -25'd13440}, '{25'd8904, 25'd7392, 25'd9072}, '{-25'd9240, 25'd10080, 25'd18816}}, '{'{-25'd10920, 25'd3696, -25'd1848}, '{25'd672, 25'd21336, 25'd11256}, '{-25'd6888, 25'd2856, -25'd8904}}, '{'{25'd3864, 25'd3360, 25'd4200}, '{25'd504, 25'd672, 25'd4032}, '{25'd4704, 25'd2184, 25'd1680}}, '{'{25'd3360, 25'd2688, 25'd1176}, '{-25'd11256, -25'd504, -25'd9912}, '{25'd336, 25'd7560, -25'd2352}}, '{'{-25'd5880, 25'd11256, 25'd1512}, '{-25'd168, 25'd9240, 25'd5880}, '{-25'd1176, 25'd6888, -25'd168}}, '{'{-25'd6048, 25'd5544, 25'd3360}, '{-25'd3528, -25'd2520, 25'd6552}, '{-25'd168, 25'd2688, 25'd504}}},
    '{'{'{-25'd7436, -25'd7175, -25'd1565}, '{-25'd8023, -25'd4762, -25'd5218}, '{-25'd4762, -25'd3848, -25'd848}}, '{'{25'd0, -25'd1696, 25'd4827}, '{25'd848, -25'd2413, -25'd2740}, '{-25'd4240, 25'd3718, 25'd1892}}, '{'{-25'd1239, -25'd130, -25'd652}, '{-25'd326, 25'd1826, -25'd4696}, '{25'd8284, -25'd4631, -25'd4827}}, '{'{-25'd6066, 25'd0, -25'd4435}, '{-25'd5675, -25'd1696, 25'd130}, '{-25'd5088, 25'd4696, -25'd5610}}, '{'{-25'd1826, -25'd4696, -25'd3066}, '{25'd2609, 25'd1239, 25'd2544}, '{-25'd3653, 25'd1370, 25'd5088}}, '{'{25'd2413, -25'd3848, -25'd4631}, '{25'd6131, -25'd4109, -25'd4762}, '{25'd1826, -25'd4044, 25'd1761}}, '{'{-25'd1305, -25'd7045, -25'd2870}, '{-25'd2022, 25'd0, -25'd4696}, '{-25'd6392, -25'd6914, -25'd4305}}, '{'{25'd717, -25'd3587, -25'd6327}, '{-25'd717, -25'd5088, 25'd522}, '{-25'd587, -25'd3131, -25'd3457}}},
    '{'{'{25'd144, -25'd13376, -25'd4027}, '{-25'd15821, -25'd6328, 25'd10931}, '{25'd3020, 25'd4602, 25'd12513}}, '{'{25'd2157, 25'd8054, 25'd2877}, '{25'd8198, 25'd2877, -25'd1870}, '{25'd7767, 25'd4027, 25'd6041}}, '{'{-25'd5178, -25'd4315, -25'd3308}, '{-25'd2014, 25'd7767, 25'd3596}, '{-25'd1151, 25'd6328, 25'd3883}}, '{'{-25'd16828, 25'd9493, -25'd431}, '{25'd14239, 25'd18266, 25'd18266}, '{-25'd11938, 25'd7911, -25'd6616}}, '{'{25'd4027, 25'd1870, 25'd575}, '{25'd7191, 25'd7479, 25'd6760}, '{25'd5753, -25'd863, 25'd4315}}, '{'{25'd6185, 25'd1438, 25'd8198}, '{-25'd6616, -25'd18410, -25'd8486}, '{25'd1438, 25'd288, -25'd3164}}, '{'{25'd863, 25'd9780, 25'd8773}, '{25'd1582, 25'd7335, -25'd719}, '{25'd3883, 25'd144, 25'd5034}}, '{'{25'd3308, -25'd575, 25'd3164}, '{25'd7048, 25'd10356, 25'd5609}, '{-25'd6185, -25'd2589, -25'd1870}}},
    '{'{'{-25'd3298, -25'd3141, 25'd9895}, '{-25'd16805, -25'd8795, 25'd14921}, '{-25'd10052, -25'd7225, -25'd15235}}, '{'{-25'd2670, 25'd2042, 25'd5968}, '{25'd471, 25'd6125, 25'd7696}, '{25'd2199, 25'd7068, -25'd2513}}, '{'{-25'd5340, 25'd5183, -25'd8481}, '{-25'd157, 25'd1571, -25'd3455}, '{-25'd2199, 25'd5497, 25'd19947}}, '{'{-25'd3455, 25'd13193, 25'd5497}, '{-25'd4869, 25'd12251, 25'd10837}, '{-25'd14607, -25'd3141, 25'd157}}, '{'{25'd6597, 25'd5811, 25'd2670}, '{25'd785, 25'd2356, 25'd4241}, '{25'd7225, 25'd1728, 25'd785}}, '{'{25'd8010, -25'd14764, 25'd1099}, '{-25'd7382, -25'd11308, -25'd1099}, '{-25'd2513, -25'd2670, -25'd8167}}, '{'{25'd1256, -25'd2670, -25'd3927}, '{25'd8481, -25'd2827, 25'd2356}, '{-25'd1099, 25'd6911, 25'd3612}}, '{'{25'd5340, 25'd5183, 25'd11622}, '{25'd15078, 25'd4555, 25'd942}, '{25'd1099, 25'd1256, 25'd3455}}},
    '{'{'{-25'd6405, -25'd1975, -25'd4190}, '{-25'd359, -25'd7543, -25'd239}, '{-25'd7662, -25'd1796, -25'd838}}, '{'{-25'd838, -25'd180, -25'd3292}, '{-25'd898, -25'd4310, 25'd60}, '{-25'd6405, 25'd1078, -25'd778}}, '{'{-25'd2394, -25'd6824, -25'd6106}, '{-25'd2215, -25'd2394, 25'd2155}, '{-25'd1556, 25'd2514, 25'd2394}}, '{'{-25'd778, -25'd1257, -25'd1197}, '{25'd658, -25'd7423, -25'd1437}, '{-25'd4729, -25'd419, -25'd2634}}, '{'{-25'd3292, -25'd4849, -25'd599}, '{25'd1796, -25'd3472, -25'd6285}, '{-25'd1796, 25'd1257, -25'd1018}}, '{'{-25'd120, -25'd5866, -25'd5028}, '{25'd838, -25'd3233, -25'd1616}, '{-25'd2813, 25'd239, 25'd1437}}, '{'{-25'd4310, -25'd5447, -25'd7483}, '{-25'd2095, 25'd1197, -25'd3472}, '{-25'd3053, 25'd658, -25'd4729}}, '{'{25'd1796, -25'd3532, 25'd1197}, '{-25'd7124, -25'd3233, -25'd6764}, '{-25'd6345, -25'd2454, -25'd4609}}},
    '{'{'{-25'd7866, 25'd2023, -25'd2397}, '{-25'd9589, -25'd7267, 25'd1873}, '{-25'd1274, 25'd300, 25'd4345}}, '{'{-25'd1199, 25'd749, 25'd2173}, '{-25'd974, -25'd4795, -25'd749}, '{25'd899, -25'd899, 25'd599}}, '{'{25'd1873, 25'd2472, 25'd2847}, '{-25'd749, 25'd3371, 25'd3446}, '{-25'd150, -25'd375, -25'd2472}}, '{'{-25'd375, 25'd2922, -25'd3596}, '{-25'd8241, 25'd4645, -25'd3671}, '{25'd1423, 25'd6068, -25'd3296}}, '{'{-25'd5244, -25'd3746, 25'd524}, '{-25'd1349, -25'd1798, -25'd6218}, '{-25'd7342, -25'd7267, -25'd3072}}, '{'{-25'd2622, -25'd2397, 25'd749}, '{-25'd5619, -25'd4570, -25'd5169}, '{-25'd974, -25'd450, -25'd6668}}, '{'{-25'd2697, 25'd0, -25'd5619}, '{-25'd3746, -25'd5019, -25'd4046}, '{-25'd5918, -25'd6743, -25'd2997}}, '{'{25'd1948, -25'd300, -25'd6143}, '{25'd3296, -25'd5844, -25'd824}, '{25'd3371, -25'd2847, -25'd1873}}},
    '{'{'{25'd834, 25'd3018, 25'd3693}, '{-25'd556, -25'd3137, 25'd2105}, '{-25'd1072, -25'd3852, 25'd3455}}, '{'{-25'd238, 25'd3217, -25'd2978}, '{-25'd2740, 25'd40, 25'd159}, '{25'd3256, -25'd3098, 25'd40}}, '{'{-25'd5083, 25'd4368, 25'd159}, '{25'd1668, 25'd3773, -25'd1271}, '{25'd3971, -25'd715, 25'd4567}}, '{'{25'd3614, -25'd4766, -25'd2780}, '{25'd437, -25'd4726, 25'd437}, '{-25'd4527, 25'd1231, -25'd2144}}, '{'{-25'd2581, -25'd1112, -25'd3971}, '{25'd3376, -25'd3574, -25'd1708}, '{-25'd1112, -25'd2899, 25'd2820}}, '{'{-25'd4408, -25'd1787, 25'd794}, '{-25'd1430, 25'd1072, -25'd1430}, '{25'd993, -25'd794, -25'd4051}}, '{'{-25'd1946, -25'd4964, -25'd2422}, '{-25'd4527, -25'd278, -25'd3852}, '{-25'd953, -25'd4527, -25'd4686}}, '{'{-25'd3614, -25'd119, -25'd40}, '{25'd3773, -25'd4090, -25'd2422}, '{25'd3733, -25'd4924, -25'd4090}}},
    '{'{'{-25'd2902, -25'd4876, -25'd2264}, '{-25'd1974, 25'd1219, -25'd1741}, '{-25'd4760, -25'd2902, -25'd3251}}, '{'{-25'd5282, -25'd6559, 25'd2032}, '{25'd0, 25'd1451, -25'd7198}, '{-25'd3018, -25'd2148, 25'd1509}}, '{'{25'd929, -25'd4644, -25'd4760}, '{-25'd7314, -25'd4412, 25'd1858}, '{-25'd639, 25'd2264, 25'd813}}, '{'{-25'd2322, -25'd406, -25'd1219}, '{-25'd6501, 25'd2438, 25'd2090}, '{-25'd3018, 25'd2496, -25'd3018}}, '{'{25'd2496, 25'd1567, -25'd1045}, '{-25'd3018, 25'd1974, -25'd4005}, '{25'd2206, 25'd522, -25'd5979}}, '{'{-25'd5631, 25'd987, 25'd987}, '{-25'd1916, -25'd7430, 25'd1858}, '{25'd1858, -25'd3599, -25'd4644}}, '{'{25'd406, -25'd813, -25'd5631}, '{-25'd1393, -25'd6792, -25'd5514}, '{-25'd4702, -25'd1335, -25'd3367}}, '{'{-25'd5224, -25'd4528, -25'd348}, '{-25'd1741, -25'd3367, -25'd871}, '{-25'd6443, -25'd1277, -25'd2380}}}
};
