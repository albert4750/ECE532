localparam bit signed [0:10][15:0] Output6 = '{-16'd31766, 16'd6828, -16'd28082, -16'd8630, 16'd2555, -16'd7124, -16'd12419, 16'd10738, -16'd4502, 16'd20481, -16'd22667};
