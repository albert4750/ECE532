localparam bit signed [0:2][0:26][19:0] Input3 = '{
    '{-20'd11, 20'd61, -20'd45, 20'd33, -20'd24, 20'd32, 20'd100, 20'd123, 20'd123, -20'd7, -20'd58, 20'd85, -20'd97, -20'd115, -20'd57, 20'd56, 20'd24, -20'd49, -20'd87, -20'd110, -20'd88, 20'd54, 20'd79, -20'd117, 20'd38, -20'd17, -20'd35},
    '{20'd121, 20'd1, 20'd95, -20'd10, -20'd84, 20'd88, -20'd3, -20'd104, -20'd61, 20'd82, 20'd111, -20'd125, 20'd106, 20'd76, 20'd102, -20'd93, 20'd86, 20'd126, 20'd61, 20'd69, 20'd87, -20'd85, -20'd96, -20'd117, -20'd24, 20'd84, 20'd10},
    '{20'd54, 20'd107, 20'd37, -20'd3, 20'd28, -20'd17, 20'd104, -20'd126, -20'd101, 20'd83, 20'd89, 20'd23, -20'd75, -20'd77, 20'd46, 20'd20, 20'd53, -20'd99, -20'd61, -20'd93, -20'd89, 20'd9, -20'd55, -20'd87, 20'd23, 20'd3, -20'd82}
};
