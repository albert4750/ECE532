logic signed [7:0] convolve17_weight[4][8][3][3] = '{
    '{
        '{'{-123, 116, -88}, '{86, 52, 43}, '{65, 6, -100}},
        '{'{5, 104, -54}, '{7, -99, -28}, '{-46, -81, 60}},
        '{'{-65, -5, 66}, '{-87, -99, -32}, '{-79, 60, -76}},
        '{'{-103, -92, 19}, '{-32, 117, -37}, '{26, -72, -72}},
        '{'{-100, 45, 87}, '{82, -123, 65}, '{-43, -94, 1}},
        '{'{-35, 109, 98}, '{-114, 106, -98}, '{9, 54, -101}},
        '{'{7, 76, -35}, '{36, 38, -36}, '{-15, -43, 87}},
        '{'{37, 20, -115}, '{-19, 40, 50}, '{105, -74, -2}}
    },
    '{
        '{'{65, -56, -70}, '{-25, -20, -55}, '{-79, -111, -79}},
        '{'{-39, 87, 57}, '{104, 121, -13}, '{74, -38, -115}},
        '{'{-97, -4, -107}, '{-31, 109, -127}, '{96, 43, 55}},
        '{'{-58, -94, 94}, '{-82, -38, 102}, '{100, 17, -16}},
        '{'{-116, -76, -81}, '{-12, 39, -16}, '{48, 55, 25}},
        '{'{-64, -68, 102}, '{30, 105, 111}, '{-28, -26, -36}},
        '{'{106, 87, -49}, '{38, -26, 86}, '{-80, -121, -91}},
        '{'{114, -62, -51}, '{-108, -82, 93}, '{-96, -76, 55}}
    },
    '{
        '{'{19, 108, 108}, '{56, -106, -42}, '{108, 101, -68}},
        '{'{34, -67, 54}, '{-90, 85, 92}, '{48, 34, 61}},
        '{'{65, 54, -19}, '{110, 17, -76}, '{-94, 43, 13}},
        '{'{-111, -97, -107}, '{98, -19, 1}, '{-59, 47, 114}},
        '{'{38, -65, 31}, '{-36, -26, 122}, '{-14, 112, -60}},
        '{'{37, 7, -61}, '{-74, -107, 21}, '{-71, 90, -62}},
        '{'{92, -81, -96}, '{101, 33, 99}, '{58, 32, -25}},
        '{'{17, 9, -29}, '{44, -42, -123}, '{86, 9, -10}}
    },
    '{
        '{'{-63, 61, 107}, '{5, 106, 68}, '{7, 54, -109}},
        '{'{114, -77, 38}, '{117, 119, 13}, '{-117, -41, -26}},
        '{'{-74, 53, -53}, '{-88, 117, -33}, '{-125, 119, 61}},
        '{'{2, 71, -126}, '{-103, -82, 5}, '{-112, -14, 8}},
        '{'{81, -8, -14}, '{-36, -50, 56}, '{-122, -51, -72}},
        '{'{92, -125, 108}, '{-69, -26, -17}, '{-124, -128, 75}},
        '{'{38, 6, -13}, '{20, 120, 70}, '{16, -64, -61}},
        '{'{-5, -59, -17}, '{-67, -89, -69}, '{80, 89, 121}}
    }
};
