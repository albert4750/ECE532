localparam bit signed [0:7][0:7][0:2][0:2][24:0] Weight2 = '{
    '{'{'{25'd3272, 25'd9452, 25'd1454}, '{-25'd11543, -25'd3908, -25'd10543}, '{-25'd4908, -25'd10816, -25'd3363}}, '{'{-25'd4635, 25'd9089, 25'd4454}, '{25'd4544, 25'd3999, -25'd1909}, '{-25'd4999, -25'd6817, -25'd5635}}, '{'{-25'd6544, 25'd182, 25'd8634}, '{25'd3545, -25'd3454, -25'd9634}, '{-25'd9907, 25'd4817, -25'd4726}}, '{'{-25'd2272, 25'd10998, -25'd5908}, '{25'd11543, 25'd8089, 25'd7453}, '{-25'd273, -25'd7998, -25'd364}}, '{'{-25'd5362, 25'd4817, 25'd1272}, '{25'd5544, 25'd6908, -25'd2545}, '{-25'd2999, -25'd1363, 25'd4363}}, '{'{-25'd2272, 25'd9362, 25'd3817}, '{25'd3999, 25'd9543, 25'd9725}, '{25'd2636, 25'd9543, 25'd9725}}, '{'{-25'd2363, -25'd3817, -25'd8907}, '{25'd9998, 25'd3999, -25'd8544}, '{25'd1182, 25'd7907, 25'd1636}}, '{'{-25'd3726, 25'd1091, 25'd91}, '{-25'd6090, 25'd3272, -25'd9634}, '{-25'd1909, 25'd2000, 25'd3545}}},
    '{'{'{25'd7125, 25'd8515, -25'd608}, '{25'd6951, 25'd8254, 25'd4866}, '{25'd608, 25'd8602, 25'd8515}}, '{'{25'd6429, -25'd8167, 25'd5300}, '{25'd2867, -25'd7993, 25'd1303}, '{25'd5821, 25'd3562, 25'd9210}}, '{'{25'd8341, -25'd782, -25'd4344}, '{25'd2520, 25'd7125, 25'd7298}, '{25'd8167, 25'd4692, 25'd7038}}, '{'{25'd11034, 25'd2520, 25'd9557}, '{-25'd1738, -25'd2607, 25'd8515}, '{25'd7993, 25'd1998, 25'd10600}}, '{'{-25'd6343, -25'd1911, 25'd261}, '{-25'd9470, -25'd1216, 25'd2867}, '{-25'd6429, 25'd1216, -25'd3562}}, '{'{25'd2085, 25'd9470, 25'd1564}, '{-25'd695, 25'd5647, -25'd2085}, '{25'd956, 25'd5821, 25'd956}}, '{'{25'd4692, 25'd7906, 25'd9905}, '{25'd10774, 25'd7298, 25'd9644}, '{-25'd3823, 25'd6603, 25'd1477}}, '{'{25'd2520, 25'd782, -25'd4431}, '{-25'd6429, -25'd695, 25'd608}, '{-25'd2433, 25'd4605, 25'd5821}}},
    '{'{'{-25'd5136, -25'd2473, -25'd3424}, '{-25'd5421, -25'd7608, 25'd4185}, '{-25'd9796, -25'd1807, -25'd9415}}, '{'{25'd8655, 25'd8084, 25'd8179}, '{-25'd9606, -25'd2473, -25'd4660}, '{25'd951, 25'd7894, 25'd4280}}, '{'{25'd7704, -25'd2568, 25'd5992}, '{25'd2283, 25'd6372, -25'd380}, '{-25'd8655, 25'd1427, 25'd4850}}, '{'{25'd0, -25'd951, -25'd2948}, '{-25'd2283, 25'd4470, 25'd2473}, '{-25'd1522, -25'd8274, 25'd666}}, '{'{25'd7799, -25'd2283, -25'd5801}, '{-25'd3614, 25'd5326, 25'd7989}, '{25'd1712, -25'd4375, 25'd5041}}, '{'{25'd3138, 25'd190, -25'd476}, '{25'd3234, 25'd761, -25'd5421}, '{-25'd6277, -25'd2948, 25'd3234}}, '{'{25'd6657, 25'd7704, -25'd4945}, '{25'd6182, 25'd7418, 25'd3234}, '{-25'd7038, -25'd12078, -25'd8559}}, '{'{-25'd285, -25'd2663, 25'd7323}, '{-25'd8179, 25'd8750, -25'd5611}, '{-25'd2853, 25'd4850, -25'd10842}}},
    '{'{'{25'd3001, -25'd4093, -25'd455}, '{-25'd4275, 25'd2729, -25'd3729}, '{25'd2638, 25'd8731, -25'd4002}}, '{'{25'd7640, 25'd7458, -25'd3456}, '{-25'd6094, -25'd3001, -25'd3365}, '{25'd3456, 25'd8095, 25'd7185}}, '{'{25'd6730, -25'd9368, 25'd5184}, '{25'd5821, -25'd9732, 25'd5002}, '{25'd2456, -25'd8368, -25'd6912}}, '{'{25'd4093, -25'd910, 25'd5821}, '{25'd3456, 25'd8004, -25'd4366}, '{25'd7276, 25'd7913, 25'd9368}}, '{'{25'd1728, 25'd5548, 25'd5548}, '{25'd3456, 25'd7185, -25'd3638}, '{25'd7640, 25'd6367, 25'd4639}}, '{'{25'd10550, 25'd6912, 25'd11096}, '{25'd3638, 25'd10369, 25'd11005}, '{25'd819, 25'd273, 25'd11551}}, '{'{25'd8731, -25'd8731, -25'd4820}, '{-25'd3183, -25'd3638, -25'd4093}, '{-25'd1910, -25'd8277, -25'd4820}}, '{'{-25'd728, 25'd4184, 25'd6185}, '{-25'd7458, 25'd5639, 25'd6185}, '{25'd9004, 25'd2092, -25'd2183}}},
    '{'{'{25'd6620, 25'd1904, 25'd725}, '{-25'd9159, -25'd5260, 25'd4444}, '{25'd5532, -25'd6711, 25'd5713}}, '{'{-25'd11608, -25'd8706, 25'd1360}, '{25'd6892, 25'd2539, -25'd272}, '{25'd4716, 25'd9431, 25'd7255}}, '{'{25'd1270, -25'd7980, -25'd1723}, '{25'd5985, 25'd3718, -25'd2539}, '{-25'd8706, 25'd7889, 25'd4444}}, '{'{-25'd3265, -25'd7799, -25'd544}, '{25'd5713, -25'd1179, 25'd7799}, '{25'd1814, 25'd6529, 25'd10338}}, '{'{-25'd4534, 25'd3627, 25'd1723}, '{-25'd6439, -25'd4897, -25'd2721}, '{25'd3899, 25'd8887, 25'd5350}}, '{'{-25'd5260, 25'd4534, -25'd10429}, '{25'd4534, 25'd4262, -25'd181}, '{-25'd8162, -25'd4625, 25'd1270}}, '{'{-25'd2086, -25'd8252, 25'd6983}, '{-25'd7255, 25'd453, 25'd5078}, '{-25'd6983, 25'd5260, 25'd6892}}, '{'{-25'd2086, -25'd9431, -25'd3083}, '{-25'd2358, 25'd6348, -25'd1814}, '{-25'd4353, 25'd544, 25'd1995}}},
    '{'{'{25'd7137, 25'd8060, 25'd8228}, '{-25'd5374, 25'd9404, 25'd4030}, '{25'd6297, 25'd3526, 25'd1343}}, '{'{25'd3778, 25'd1595, -25'd2603}, '{25'd9320, 25'd3694, 25'd7053}, '{-25'd5709, -25'd4954, 25'd9320}}, '{'{25'd1427, 25'd5709, -25'd10747}, '{25'd3694, 25'd6297, 25'd4198}, '{-25'd6885, -25'd5122, 25'd4366}}, '{'{25'd168, 25'd4030, -25'd2435}, '{25'd9236, 25'd9320, 25'd8312}, '{25'd7389, -25'd672, 25'd9740}}, '{'{-25'd1343, -25'd7809, 25'd10243}, '{25'd252, 25'd3526, -25'd6213}, '{25'd6297, 25'd8396, -25'd7725}}, '{'{25'd9992, 25'd10160, 25'd10160}, '{25'd9992, 25'd5961, 25'd6549}, '{25'd10160, 25'd10411, 25'd3359}}, '{'{-25'd5458, 25'd5206, 25'd5877}, '{25'd1427, -25'd6465, -25'd4450}, '{-25'd1763, 25'd9824, 25'd1427}}, '{'{-25'd5626, -25'd5122, -25'd6969}, '{25'd3191, 25'd9824, -25'd5626}, '{-25'd6297, -25'd3107, 25'd2099}}},
    '{'{'{25'd7835, 25'd5252, 25'd8437}, '{25'd1722, -25'd3099, 25'd2411}, '{25'd1636, 25'd1291, -25'd4649}}, '{'{25'd5768, 25'd1291, -25'd3960}, '{25'd3530, 25'd172, -25'd7318}, '{25'd4477, -25'd7490, 25'd1033}}, '{'{-25'd3702, 25'd1636, -25'd430}, '{25'd1378, 25'd1464, -25'd10590}, '{25'd6113, -25'd5768, -25'd1808}}, '{'{25'd7662, 25'd6113, 25'd7060}, '{25'd3788, -25'd4391, 25'd861}, '{25'd1808, -25'd2238, -25'd861}}, '{'{25'd1636, -25'd4994, -25'd1636}, '{-25'd8954, -25'd3358, 25'd8179}, '{25'd9643, -25'd4994, 25'd5941}}, '{'{25'd8265, -25'd3099, 25'd9298}, '{25'd8782, 25'd9212, -25'd603}, '{25'd4133, 25'd2669, 25'd10934}}, '{'{-25'd775, 25'd2325, -25'd344}, '{25'd4735, 25'd3702, 25'd7404}, '{25'd775, -25'd9126, 25'd0}}, '{'{25'd6888, -25'd6974, -25'd4821}, '{25'd7490, -25'd2755, -25'd86}, '{-25'd603, 25'd7060, 25'd4391}}},
    '{'{'{-25'd2108, 25'd2186, -25'd7103}, '{-25'd2264, -25'd9211, -25'd2498}, '{-25'd8352, -25'd9367, -25'd2966}}, '{'{25'd9913, 25'd6166, -25'd7493}, '{-25'd6635, 25'd2810, -25'd5230}, '{-25'd6713, -25'd1093, -25'd6947}}, '{'{-25'd3825, -25'd5854, -25'd4996}, '{25'd7181, 25'd1015, 25'd1483}, '{-25'd6166, -25'd9913, 25'd1717}}, '{'{-25'd4839, 25'd624, -25'd7337}, '{-25'd2342, -25'd5698, 25'd6869}, '{-25'd8040, -25'd7259, -25'd6401}}, '{'{-25'd9367, -25'd8196, 25'd8196}, '{25'd8586, 25'd6947, -25'd9757}, '{-25'd3903, 25'd8586, -25'd78}}, '{'{-25'd2966, -25'd9913, 25'd3825}, '{25'd2029, -25'd4215, -25'd2342}, '{25'd1873, 25'd1561, -25'd6323}}, '{'{25'd4527, 25'd6713, 25'd1873}, '{-25'd6010, 25'd1405, -25'd2264}, '{25'd937, 25'd1873, -25'd4683}}, '{'{25'd3903, 25'd9133, -25'd156}, '{-25'd7493, -25'd3591, 25'd1873}, '{-25'd3747, 25'd1795, 25'd2576}}}
};
