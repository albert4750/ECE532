`ifndef ECE532_CONSTANTS_SVH
`define ECE532_CONSTANTS_SVH

package constants;

    parameter int DSPInAWidth = 25;
    parameter int DSPInBWidth = 18;
    parameter int DSPOutWidth = 48;

endpackage : constants

`endif  // ECE532_CONSTANTS_SVH
