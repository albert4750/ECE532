localparam bit signed [0:15][7:0] Output8 = '{40, -101, 86, -110, 100, 24, -37, 95, -117, 47, 113, 109, -60, 61, 24, -59};
