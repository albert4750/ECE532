localparam bit signed [0:63][47:0] Bias1 = '{48'd166226, -48'd183914, -48'd56920, -48'd53351, 48'd90429, 48'd175172, 48'd57623, 48'd186039, -48'd175720, -48'd190112, -48'd105777, -48'd188342, 48'd154547, 48'd182465, 48'd125648, 48'd167798, 48'd55580, 48'd121001, -48'd180550, 48'd168617, -48'd137409, 48'd3929, 48'd56941, -48'd181172, 48'd139485, -48'd127733, -48'd160746, 48'd157616, -48'd142582, 48'd177469, 48'd167471, -48'd2743, 48'd180717, 48'd75439, -48'd47180, -48'd110262, 48'd36936, -48'd8294, -48'd155427, -48'd185096, -48'd150926, 48'd102696, 48'd28220, 48'd93235, -48'd159354, 48'd155794, 48'd174163, 48'd104811, 48'd133538, -48'd168175, 48'd89507, -48'd9392, -48'd168361, -48'd163505, 48'd57009, -48'd133867, 48'd66084, 48'd40202, -48'd20299, -48'd179926, -48'd163776, 48'd109338, 48'd101394, -48'd122617};
