localparam bit signed [0:2][0:26][19:0] Input4 = '{
    '{20'd90, 20'd50, -20'd20, -20'd125, -20'd97, -20'd119, 20'd10, -20'd101, 20'd45, 20'd71, 20'd39, -20'd67, -20'd43, -20'd31, -20'd84, -20'd94, 20'd34, -20'd40, -20'd95, 20'd5, 20'd104, 20'd127, -20'd92, -20'd128, 20'd75, -20'd94, 20'd69},
    '{-20'd2, 20'd53, 20'd126, -20'd48, 20'd62, 20'd8, 20'd61, 20'd1, 20'd81, -20'd16, -20'd93, -20'd8, -20'd37, 20'd40, -20'd12, -20'd92, 20'd48, -20'd103, -20'd61, -20'd25, 20'd124, -20'd93, -20'd14, -20'd98, -20'd99, 20'd113, -20'd95},
    '{20'd18, -20'd111, 20'd93, -20'd44, 20'd125, -20'd126, -20'd59, -20'd27, 20'd12, -20'd84, -20'd11, 20'd125, -20'd62, -20'd17, -20'd37, -20'd43, 20'd39, -20'd89, 20'd75, 20'd22, 20'd30, 20'd17, 20'd70, 20'd71, -20'd110, -20'd36, -20'd85}
};
