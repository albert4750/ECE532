localparam bit signed [0:26][19:0] Output6 = '{-20'd267, 20'd143, 20'd146, 20'd171, 20'd47, 20'd95, -20'd42, -20'd116, -20'd10, -20'd192, -20'd83, 20'd46, -20'd109, -20'd284, 20'd54, 20'd43, -20'd70, 20'd203, -20'd201, 20'd51, 20'd104, -20'd149, 20'd31, 20'd30, 20'd71, -20'd177, 20'd92};
