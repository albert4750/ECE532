localparam bit signed [0:146][7:0] Input9 = '{-31, 14, -122, -40, 118, -125, -60, -27, 104, -33, 27, -14, 105, -61, -94, 41, -115, -1, -15, 17, -22, 40, 109, 74, -90, -86, -61, -101, 60, 15, 114, 34, 100, 106, -25, 50, -84, -44, -76, 25, 75, 44, -47, 127, 5, -45, 71, 127, -60, -33, -35, -22, 114, -37, 32, 107, 41, 82, 29, 13, 114, -20, 9, -74, 8, -103, 33, -111, 113, 47, -112, -79, -66, -57, -34, 126, 80, -42, 123, 37, -119, 46, 12, -40, -3, -11, 22, 56, -50, -83, -95, 62, -124, -59, -3, -52, 41, 12, -128, 69, 22, 105, -31, 49, -13, -63, 10, 70, -6, -112, 71, 27, -90, -21, -44, 41, 82, -13, 106, 70, 38, 34, -15, 74, 127, -25, -88, -88, 27, -34, 123, 36, -30, -69, -39, 27, 56, -1, 58, -97, -80, 107, -2, 3, -64, -91, 119};
