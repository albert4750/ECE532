logic signed [7:0] convolve8_weight[4][8][3][3] = '{
    '{
        '{'{91, 103, -30}, '{-57, -34, -83}, '{80, -63, -40}},
        '{'{-112, -83, -1}, '{91, 37, 50}, '{24, 48, 76}},
        '{'{-124, 112, 51}, '{46, -88, 14}, '{113, 10, 27}},
        '{'{-50, -26, 13}, '{-124, 86, -113}, '{-99, 78, 42}},
        '{'{25, 75, 95}, '{91, -106, -18}, '{-85, 84, 55}},
        '{'{125, 2, 25}, '{-3, -8, 0}, '{-33, 56, -18}},
        '{'{70, 82, -42}, '{62, 127, -82}, '{123, -39, 77}},
        '{'{12, -66, -91}, '{83, 31, -9}, '{28, -69, 120}}
    },
    '{
        '{'{-45, -88, -24}, '{-7, -39, 111}, '{-99, -100, -76}},
        '{'{-86, 10, 84}, '{-111, 0, 39}, '{-90, 98, 65}},
        '{'{-80, 86, -83}, '{-6, 49, -106}, '{103, 126, -36}},
        '{'{-63, -43, -62}, '{-96, 50, -58}, '{-26, 35, 117}},
        '{'{100, 23, 115}, '{-6, -46, -26}, '{-39, 110, -49}},
        '{'{-15, 27, -43}, '{-127, -119, -13}, '{-47, 11, -64}},
        '{'{119, -61, 121}, '{61, -74, -92}, '{84, -2, -109}},
        '{'{111, 69, 84}, '{-3, 62, 68}, '{41, 80, 16}}
    },
    '{
        '{'{57, 5, -32}, '{-106, 3, 8}, '{-66, -36, 41}},
        '{'{-54, -26, -36}, '{-33, -20, 11}, '{34, -37, -79}},
        '{'{-57, 39, -26}, '{-9, -70, -123}, '{-55, -40, 12}},
        '{'{104, 97, -69}, '{78, 109, -113}, '{-124, 22, 52}},
        '{'{-62, -57, -19}, '{-56, -123, -89}, '{-49, -49, -87}},
        '{'{89, 22, 89}, '{89, 19, -66}, '{-99, -119, 11}},
        '{'{-3, -29, -102}, '{-25, 127, 82}, '{-56, 127, 1}},
        '{'{-29, -14, 113}, '{46, -73, -118}, '{74, -104, 127}}
    },
    '{
        '{'{-33, -85, 91}, '{13, 78, -73}, '{-123, 23, -86}},
        '{'{-25, -79, -27}, '{-26, -53, -11}, '{56, 43, 24}},
        '{'{-47, -107, 94}, '{18, -65, -39}, '{-99, -91, 49}},
        '{'{40, 113, -22}, '{95, -25, -117}, '{-72, 117, 63}},
        '{'{14, -96, 65}, '{-7, -11, -63}, '{-92, 122, -103}},
        '{'{76, -56, -78}, '{-116, 24, 19}, '{67, 10, -121}},
        '{'{52, -36, -114}, '{72, -82, 99}, '{-93, 81, 23}},
        '{'{-67, -11, 53}, '{-116, 45, -121}, '{122, 47, -18}}
    }
};
