wire signed [7:0] convolve2_weight[4][8][3][3];
assign convolve2_weight = '{'{'{'{75, 22, 30}, '{17, 70, 71}, '{-110, -36, -85}}, '{'{-45, 49, -87}, '{-35, 46, 21}, '{73, -39, 114}}, '{'{96, 91, -55}, '{-100, 107, 81}, '{-23, 58, 0}}, '{'{86, -65, -112}, '{-22, 36, -34}, '{-104, -12, 63}}, '{'{67, -77, 8}, '{56, -37, -35}, '{-5, 110, -41}}, '{'{32, 19, -56}, '{71, -41, -115}, '{-70, -47, -8}}, '{'{-12, 55, -64}, '{75, 92, 36}, '{-103, -96, 42}}, '{'{-114, 86, -100}, '{-108, 82, -60}, '{-106, 99, -6}}}, '{'{'{-45, 7, 72}, '{-67, 13, -123}, '{-128, 8, 79}}, '{'{79, 53, 11}, '{-124, 39, -36}, '{45, -102, -54}}, '{'{-76, 110, 49}, '{91, -77, 99}, '{-23, -110, -11}}, '{'{-94, -77, 30}, '{53, -70, 43}, '{-73, 124, 124}}, '{'{-110, 45, -41}, '{65, -58, 106}, '{-75, -80, -34}}, '{'{-69, -48, 26}, '{-4, 35, -70}, '{49, -22, 73}}, '{'{-84, -115, -7}, '{-58, -90, 39}, '{8, -115, 120}}, '{'{7, 80, 120}, '{-106, 120, -49}, '{89, -120, 99}}}, '{'{'{-122, 81, 71}, '{84, 89, 66}, '{-68, 16, -72}}, '{'{-14, 109, 23}, '{-104, -124, -28}, '{108, -79, -41}}, '{'{-98, -74, 25}, '{-108, -31, -27}, '{57, 23, 27}}, '{'{-99, 33, -13}, '{-75, -9, 51}, '{-42, 118, -121}}, '{'{-23, 113, 9}, '{54, 0, -45}, '{-8, 36, 81}}, '{'{20, -11, 112}, '{-125, -2, -86}, '{-63, -108, -92}}, '{'{-60, 80, -16}, '{47, 10, 109}, '{-24, 94, -37}}, '{'{-85, -65, 31}, '{20, 70, -119}, '{60, -37, -17}}}, '{'{'{35, -45, -52}, '{-110, -15, -54}, '{98, 97, 43}}, '{'{3, 12, 100}, '{-70, 1, -15}, '{0, -89, -104}}, '{'{58, -92, -29}, '{-59, 6, -125}, '{98, -7, 40}}, '{'{60, 33, -100}, '{-60, -102, 96}, '{120, -19, 51}}, '{'{73, 53, 69}, '{33, 7, -3}, '{-34, -56, 118}}, '{'{-44, 7, 67}, '{85, 91, -20}, '{-61, -26, -44}}, '{'{-57, -45, 95}, '{-128, 5, -37}, '{-21, 30, 73}}, '{'{83, -121, 21}, '{101, 92, 8}, '{43, -82, -128}}}};
