logic signed [15:0] layer2_weight[8][16][1][1] = '{
    '{
        '{'{-3226}},
        '{'{26187}},
        '{'{-14475}},
        '{'{23480}},
        '{'{32171}},
        '{'{-28520}},
        '{'{-12975}},
        '{'{30229}},
        '{'{-10274}},
        '{'{19602}},
        '{'{12351}},
        '{'{21849}},
        '{'{1565}},
        '{'{-8923}},
        '{'{-13391}},
        '{'{-11096}}
    },
    '{
        '{'{-28175}},
        '{'{-22166}},
        '{'{23775}},
        '{'{20583}},
        '{'{3339}},
        '{'{24888}},
        '{'{24565}},
        '{'{7615}},
        '{'{22670}},
        '{'{-23264}},
        '{'{6337}},
        '{'{-27527}},
        '{'{-16011}},
        '{'{-31935}},
        '{'{22564}},
        '{'{-18694}}
    },
    '{
        '{'{-30695}},
        '{'{-20532}},
        '{'{-26552}},
        '{'{30770}},
        '{'{14860}},
        '{'{2968}},
        '{'{12435}},
        '{'{-2365}},
        '{'{-9846}},
        '{'{-9721}},
        '{'{-15436}},
        '{'{-17316}},
        '{'{-498}},
        '{'{-13880}},
        '{'{-4050}},
        '{'{5347}}
    },
    '{
        '{'{12323}},
        '{'{2257}},
        '{'{-31593}},
        '{'{10301}},
        '{'{-10635}},
        '{'{17589}},
        '{'{-11764}},
        '{'{5549}},
        '{'{32263}},
        '{'{29178}},
        '{'{-10833}},
        '{'{-22418}},
        '{'{-7513}},
        '{'{32606}},
        '{'{5779}},
        '{'{1258}}
    },
    '{
        '{'{1901}},
        '{'{-27726}},
        '{'{-16831}},
        '{'{19371}},
        '{'{16978}},
        '{'{-14898}},
        '{'{30715}},
        '{'{-2983}},
        '{'{101}},
        '{'{-5768}},
        '{'{20664}},
        '{'{-17848}},
        '{'{6834}},
        '{'{10274}},
        '{'{17370}},
        '{'{8715}}
    },
    '{
        '{'{-13716}},
        '{'{3211}},
        '{'{-22168}},
        '{'{6564}},
        '{'{-12418}},
        '{'{19633}},
        '{'{-12340}},
        '{'{22481}},
        '{'{21727}},
        '{'{20426}},
        '{'{5936}},
        '{'{-11702}},
        '{'{-4981}},
        '{'{-17827}},
        '{'{5666}},
        '{'{13002}}
    },
    '{
        '{'{3532}},
        '{'{2801}},
        '{'{-25305}},
        '{'{26992}},
        '{'{-6646}},
        '{'{25346}},
        '{'{-6791}},
        '{'{-27665}},
        '{'{75}},
        '{'{-30802}},
        '{'{19507}},
        '{'{23028}},
        '{'{12201}},
        '{'{-28678}},
        '{'{31835}},
        '{'{3715}}
    },
    '{
        '{'{18704}},
        '{'{-17089}},
        '{'{-17600}},
        '{'{7949}},
        '{'{-28890}},
        '{'{-28412}},
        '{'{-17917}},
        '{'{25491}},
        '{'{21073}},
        '{'{-29552}},
        '{'{-30338}},
        '{'{31559}},
        '{'{8856}},
        '{'{9483}},
        '{'{-8042}},
        '{'{-12740}}
    }
};
