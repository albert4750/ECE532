localparam bit signed [0:26][19:0] Output2 = '{-20'd3, -20'd76, 20'd149, -20'd86, -20'd173, 20'd70, 20'd35, 20'd191, 20'd139, -20'd165, 20'd47, -20'd159, -20'd136, -20'd202, 20'd12, -20'd47, -20'd83, -20'd269, -20'd77, -20'd83, -20'd152, -20'd253, -20'd213, -20'd24, -20'd10, 20'd113, 20'd110};
