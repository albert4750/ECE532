logic signed [7:0] convolve15_weight[4][8][3][3] = '{
    '{
        '{'{105, 5, 88}, '{127, -45, 54}, '{101, -125, -45}},
        '{'{23, -80, -34}, '{30, 89, 7}, '{42, 12, -124}},
        '{'{112, 27, 76}, '{-17, 74, 124}, '{43, 53, 110}},
        '{'{10, 115, -85}, '{-122, 71, -128}, '{-77, 34, -32}},
        '{'{-105, 64, 71}, '{30, -110, -96}, '{-126, 38, -116}},
        '{'{-64, -2, 124}, '{-56, -125, 13}, '{-2, 90, 3}},
        '{'{102, 70, 6}, '{20, -70, -126}, '{85, 47, 127}},
        '{'{52, -70, -18}, '{-46, 126, -48}, '{-71, 43, -95}}
    },
    '{
        '{'{106, -59, 93}, '{-49, -39, 109}, '{117, -104, -28}},
        '{'{60, -7, -64}, '{61, -51, -116}, '{70, -15, -79}},
        '{'{3, 32, -13}, '{49, 99, 13}, '{-53, -111, -60}},
        '{'{87, -81, -54}, '{38, -12, 117}, '{-26, 48, -92}},
        '{'{93, -103, -93}, '{71, 64, -64}, '{-120, 67, -122}},
        '{'{-27, 124, 7}, '{51, 77, -46}, '{-8, -111, -125}},
        '{'{-2, -120, -81}, '{-85, 61, -125}, '{-84, -53, 117}},
        '{'{-79, -78, 10}, '{43, 79, 91}, '{-26, -66, 99}}
    },
    '{
        '{'{-46, 125, -66}, '{-11, 35, -43}, '{28, 59, 97}},
        '{'{-39, 74, -127}, '{122, 21, 25}, '{10, -8, 41}},
        '{'{-115, 51, -62}, '{82, 84, 7}, '{-88, -72, -43}},
        '{'{-91, 46, 83}, '{90, 55, 6}, '{-128, 8, 124}},
        '{'{85, -5, 111}, '{37, 67, 46}, '{104, 41, -36}},
        '{'{-65, -71, 119}, '{-28, -89, 65}, '{51, 61, -19}},
        '{'{69, 58, -37}, '{-33, 40, -55}, '{53, -8, -121}},
        '{'{-29, 47, 69}, '{41, -100, 118}, '{-6, -43, -117}}
    },
    '{
        '{'{-125, -110, 35}, '{-82, -23, 17}, '{-17, 27, -74}},
        '{'{-17, 73, 19}, '{71, -57, -27}, '{43, 126, 44}},
        '{'{-18, 46, 34}, '{33, -54, -9}, '{-59, 92, -82}},
        '{'{32, 83, 39}, '{30, 95, -17}, '{47, 1, 32}},
        '{'{-2, -24, -15}, '{63, -9, -83}, '{55, -18, -10}},
        '{'{-64, -27, 85}, '{22, 27, -123}, '{-19, -93, -19}},
        '{'{-93, -4, -24}, '{67, 28, -37}, '{123, 9, -85}},
        '{'{3, -21, 11}, '{51, 86, -22}, '{106, 4, 29}}
    }
};
