localparam bit signed [0:63][0:2][0:8][0:8][24:0] Weight1 = '{
    '{'{'{25'd915352, 25'd1464563, -25'd3075583, 25'd3148811, 25'd4430304, -25'd439369, 25'd3624794, 25'd3405109, 25'd622439}, '{-25'd2306687, -25'd3038969, 25'd1391335, 25'd1391335, 25'd439369, 25'd4283847, -25'd842124, -25'd3917706, 25'd1940546}, '{-25'd878738, -25'd2929126, 25'd1830704, -25'd878738, -25'd3624794, -25'd2123617, 25'd3954321, 25'd4064163, 25'd3331881}, '{25'd2087002, 25'd1391335, 25'd1208265, -25'd146456, 25'd3917706, -25'd1135036, -25'd2526371, -25'd439369, 25'd2929126}, '{25'd915352, 25'd4283847, 25'd1940546, 25'd3368495, 25'd4100777, -25'd2672828, 25'd2819284, 25'd1647634, 25'd1574405}, '{25'd2562986, 25'd439369, -25'd512597, -25'd768896, 25'd3661408, -25'd2306687, -25'd329527, 25'd3368495, 25'd1757476}, '{-25'd1830704, -25'd549211, 25'd2892512, -25'd1903932, 25'd4247233, 25'd3807864, 25'd549211, 25'd3661408, 25'd2526371}, '{-25'd1244879, 25'd4100777, -25'd951966, 25'd1208265, -25'd1611019, 25'd2636214, -25'd1830704, -25'd2270073, -25'd585825}, '{-25'd1720862, -25'd549211, 25'd805510, 25'd2636214, -25'd585825, -25'd3112197, -25'd585825, 25'd3405109, -25'd3368495}}, '{'{25'd366141, 25'd842124, 25'd622439, -25'd2929126, 25'd2489757, -25'd1354721, 25'd3038969, -25'd439369, 25'd2013774}, '{25'd1061808, -25'd475983, -25'd3478337, 25'd1098422, -25'd2709442, 25'd2562986, 25'd3954321, 25'd2599600, 25'd439369}, '{-25'd366141, -25'd659053, 25'd4357075, 25'd3807864, -25'd2087002, -25'd1135036, -25'd402755, -25'd3441723, 25'd3148811}, '{-25'd3222039, -25'd622439, 25'd146456, 25'd3990935, -25'd1867318, 25'd2636214, -25'd3185425, 25'd3295267, -25'd2929126}, '{-25'd2709442, -25'd1354721, 25'd402755, 25'd951966, 25'd1464563, -25'd1611019, 25'd1427949, 25'd146456, 25'd1977160}, '{-25'd2343301, -25'd3624794, -25'd3954321, 25'd4540146, -25'd3222039, -25'd2050388, 25'd3551566, -25'd1025194, -25'd2929126}, '{-25'd3258653, 25'd256299, 25'd3807864, 25'd109842, 25'd4503532, -25'd3771250, 25'd1537791, 25'd4064163, -25'd512597}, '{-25'd3990935, -25'd1537791, 25'd3002354, -25'd549211, 25'd1684248, -25'd1647634, 25'd329527, -25'd329527, -25'd3771250}, '{25'd2123617, 25'd3405109, -25'd109842, 25'd3990935, -25'd3405109, 25'd4174005, 25'd1061808, -25'd659053, -25'd1098422}}, '{'{25'd1098422, 25'd1684248, 25'd1098422, -25'd915352, 25'd3624794, 25'd3551566, 25'd1098422, -25'd3038969, -25'd1830704}, '{-25'd402755, -25'd402755, -25'd1830704, 25'd3258653, 25'd1391335, -25'd3038969, 25'd1574405, -25'd2416529, 25'd951966}, '{25'd3954321, -25'd878738, 25'd3295267, 25'd3588180, 25'd2453143, 25'd2599600, 25'd219684, 25'd951966, -25'd3734636}, '{-25'd3917706, -25'd475983, -25'd2746056, 25'd1391335, 25'd951966, -25'd2416529, -25'd1574405, 25'd2087002, 25'd3075583}, '{25'd3441723, 25'd1354721, 25'd805510, -25'd842124, 25'd878738, -25'd622439, -25'd3368495, -25'd146456, 25'd36614}, '{25'd585825, 25'd402755, -25'd219684, 25'd4649988, 25'd1427949, 25'd3038969, 25'd0, -25'd1244879, -25'd2526371}, '{25'd2965740, 25'd2196845, 25'd73228, 25'd329527, 25'd2160231, 25'd3514952, 25'd1391335, -25'd2343301, -25'd1611019}, '{-25'd3478337, 25'd1684248, -25'd366141, 25'd1501177, -25'd3624794, -25'd768896, 25'd2013774, 25'd2636214, 25'd3112197}, '{-25'd2306687, -25'd1611019, 25'd878738, 25'd3954321, -25'd146456, -25'd1611019, 25'd292913, -25'd256299, -25'd2965740}}},
    '{'{'{-25'd3724829, -25'd3925089, -25'd3564621, 25'd3925089, -25'd2242908, 25'd2443167, 25'd4045244, -25'd3724829, 25'd720935}, '{-25'd1441869, 25'd3164102, 25'd1001298, -25'd160208, 25'd1041350, -25'd2603375, 25'd3364362, -25'd2643427, 25'd2282960}, '{25'd1762285, -25'd1682181, -25'd1121454, 25'd1481921, 25'd4005192, -25'd2162804, -25'd3043946, -25'd760987, -25'd2122752}, '{25'd2042648, -25'd2723531, 25'd1161506, 25'd1562025, -25'd3244206, -25'd1882440, -25'd1802337, -25'd760987, 25'd120156}, '{25'd720935, 25'd2843687, -25'd2202856, 25'd120156, 25'd1361765, 25'd881142, 25'd1602077, -25'd3164102, 25'd4165400}, '{25'd4245504, 25'd2403115, -25'd3684777, 25'd4605971, -25'd3244206, -25'd2603375, -25'd881142, 25'd1521973, 25'd3724829}, '{25'd1161506, -25'd720935, -25'd1842388, 25'd2042648, -25'd2002596, -25'd1562025, -25'd40052, 25'd2843687, -25'd1081402}, '{-25'd1762285, -25'd1962544, 25'd2683479, -25'd1682181, 25'd921194, -25'd1722233, 25'd2643427, -25'd3404414, -25'd1562025}, '{25'd1642129, -25'd1401817, 25'd2082700, 25'd2803635, 25'd1401817, -25'd2723531, 25'd2963842, 25'd4445764, 25'd3284258}}, '{'{25'd2042648, -25'd1441869, -25'd3364362, -25'd2363063, 25'd1842388, -25'd80104, -25'd2483219, 25'd3925089, -25'd2683479}, '{-25'd440571, 25'd4085296, 25'd760987, 25'd2002596, 25'd3164102, 25'd2122752, 25'd2323012, -25'd2603375, -25'd2643427}, '{25'd4085296, 25'd2122752, -25'd1802337, 25'd3244206, 25'd440571, -25'd2843687, 25'd2162804, -25'd3164102, 25'd3164102}, '{25'd2002596, 25'd3124050, -25'd2242908, 25'd4605971, 25'd3925089, 25'd2282960, 25'd4605971, -25'd2563323, -25'd1121454}, '{25'd4245504, 25'd4245504, -25'd1842388, 25'd4806231, -25'd1962544, 25'd2042648, 25'd1281662, -25'd2042648, -25'd1802337}, '{-25'd3844985, 25'd1401817, 25'd5046542, 25'd2162804, 25'd320415, 25'd1281662, 25'd5006490, 25'd2563323, -25'd2443167}, '{-25'd1682181, 25'd1802337, 25'd1161506, -25'd1682181, -25'd2443167, 25'd2763583, 25'd3844985, -25'd1602077, 25'd801038}, '{-25'd1361765, 25'd2202856, 25'd600779, 25'd2282960, -25'd2923790, -25'd2162804, 25'd680883, 25'd961246, -25'd3164102}, '{-25'd80104, -25'd3444465, -25'd680883, -25'd3644725, -25'd2643427, -25'd560727, 25'd1361765, -25'd4165400, 25'd480623}}, '{'{25'd2323012, 25'd3764881, -25'd3965140, -25'd3284258, 25'd3444465, 25'd2082700, 25'd1201558, 25'd3404414, -25'd3965140}, '{-25'd1962544, 25'd1802337, 25'd3043946, -25'd4245504, -25'd3524569, 25'd3885037, 25'd1682181, -25'd1642129, 25'd2122752}, '{25'd2563323, 25'd440571, 25'd280363, 25'd2122752, 25'd1401817, -25'd2923790, 25'd720935, 25'd1081402, -25'd4285556}, '{25'd1602077, 25'd1161506, 25'd320415, -25'd2323012, -25'd2763583, 25'd2242908, 25'd1001298, 25'd160208, -25'd3804933}, '{-25'd3564621, 25'd2363063, 25'd120156, 25'd1201558, 25'd2643427, 25'd1201558, -25'd2483219, -25'd720935, 25'd2363063}, '{-25'd3965140, 25'd3684777, 25'd3364362, -25'd2242908, -25'd2242908, 25'd4646023, 25'd3644725, -25'd2122752, -25'd801038}, '{-25'd1922492, -25'd1802337, -25'd1201558, 25'd1121454, 25'd680883, 25'd841090, 25'd2403115, -25'd2643427, -25'd480623}, '{-25'd3965140, -25'd3564621, 25'd1562025, -25'd3124050, -25'd3043946, 25'd480623, -25'd1161506, -25'd3244206, -25'd5086594}, '{25'd3885037, 25'd560727, -25'd4085296, 25'd2723531, -25'd4125348, 25'd1802337, 25'd2643427, 25'd1762285, -25'd3164102}}},
    '{'{'{25'd2257358, -25'd3103867, 25'd451472, -25'd1918754, 25'd2257358, -25'd2652395, -25'd1580150, 25'd1467282, -25'd3386036}, '{-25'd3724640, 25'd3611772, 25'd3781074, 25'd2652395, 25'd3329602, 25'd3160301, 25'd2652395, 25'd451472, -25'd2483093}, '{-25'd2144490, 25'd507905, 25'd1749452, -25'd1128679, 25'd2088056, -25'd1975188, -25'd2990999, 25'd2483093, 25'd620773}, '{25'd2426659, 25'd395038, 25'd2370225, -25'd1185113, -25'd790075, -25'd1862320, -25'd4345413, 25'd282170, -25'd2934565}, '{25'd3160301, -25'd3216735, 25'd0, 25'd3329602, 25'd4909753, -25'd790075, 25'd2370225, -25'd1523716, -25'd4796885}, '{25'd2483093, -25'd56434, 25'd1523716, 25'd1805886, 25'd3555338, 25'd620773, 25'd2652395, -25'd1467282, -25'd4288979}, '{-25'd4966187, 25'd959377, 25'd3724640, 25'd1918754, -25'd959377, 25'd3103867, 25'd3273168, 25'd1805886, -25'd3103867}, '{-25'd3047433, -25'd677207, -25'd1749452, 25'd620773, 25'd2652395, 25'd3103867, -25'd2257358, 25'd2708829, -25'd2765263}, '{25'd2370225, -25'd112868, 25'd2708829, -25'd2765263, 25'd4288979, 25'd2483093, -25'd2257358, -25'd4063244, 25'd2765263}}, '{'{25'd1072245, -25'd1975188, -25'd2257358, -25'd3103867, -25'd2652395, 25'd3273168, 25'd1185113, 25'd677207, 25'd2539527}, '{25'd3386036, -25'd2539527, -25'd395038, 25'd1467282, 25'd5643394, 25'd564339, -25'd564339, -25'd2878131, -25'd4571149}, '{25'd1749452, 25'd2370225, -25'd3216735, 25'd4571149, 25'd5079055, -25'd2878131, -25'd2539527, 25'd451472, -25'd733641}, '{-25'd1636584, 25'd3555338, 25'd4571149, 25'd2539527, 25'd2031622, -25'd1297981, 25'd1805886, -25'd2990999, -25'd3668206}, '{-25'd338604, -25'd3047433, 25'd3893942, 25'd3950376, 25'd5812696, 25'd5756262, 25'd56434, 25'd3724640, -25'd902943}, '{25'd1918754, -25'd1636584, -25'd2934565, 25'd2426659, 25'd2539527, -25'd225736, -25'd2539527, -25'd5135488, -25'd2200924}, '{25'd1693018, 25'd1467282, 25'd4514715, 25'd4401847, 25'd2765263, -25'd1128679, -25'd395038, -25'd1297981, -25'd3724640}, '{25'd846509, -25'd2652395, 25'd0, -25'd2765263, -25'd1975188, -25'd564339, 25'd1749452, -25'd4345413, 25'd169302}, '{-25'd1072245, 25'd1128679, 25'd846509, 25'd1862320, 25'd2765263, 25'd3103867, -25'd4119678, -25'd2934565, -25'd2765263}}, '{'{-25'd1297981, 25'd395038, -25'd1580150, -25'd1862320, 25'd6094865, 25'd3668206, -25'd3442470, -25'd451472, -25'd3273168}, '{25'd282170, -25'd2708829, -25'd3160301, -25'd902943, 25'd2483093, 25'd5022621, 25'd225736, -25'd2370225, -25'd1241547}, '{25'd3216735, 25'd1523716, -25'd1467282, 25'd6320601, 25'd3498904, -25'd564339, 25'd1693018, -25'd2257358, -25'd733641}, '{25'd1749452, -25'd733641, 25'd4401847, 25'd5925564, 25'd4401847, 25'd2370225, 25'd2426659, -25'd1975188, -25'd2878131}, '{-25'd3668206, -25'd169302, -25'd1467282, 25'd4401847, 25'd2652395, -25'd282170, 25'd6546337, 25'd1523716, -25'd2313792}, '{-25'd3498904, 25'd1354415, -25'd1523716, 25'd7167110, 25'd2200924, 25'd3103867, -25'd1580150, -25'd1749452, -25'd3047433}, '{25'd3442470, -25'd225736, -25'd1241547, 25'd5586960, 25'd733641, -25'd1410848, -25'd1862320, -25'd4288979, -25'd3273168}, '{-25'd1467282, -25'd225736, 25'd3781074, -25'd959377, 25'd620773, 25'd338604, -25'd3498904, -25'd4684017, -25'd1805886}, '{-25'd1410848, 25'd3216735, -25'd225736, -25'd2652395, 25'd3047433, 25'd507905, 25'd4119678, -25'd5417658, 25'd2031622}}},
    '{'{'{25'd3808688, 25'd754551, 25'd1832482, 25'd2012137, 25'd3880550, 25'd3629033, -25'd718620, 25'd826414, 25'd2946344}, '{25'd1652827, 25'd431172, 25'd3305654, 25'd2012137, 25'd4491378, -25'd2838551, 25'd1113862, 25'd1868413, -25'd503034}, '{-25'd1473172, 25'd467103, 25'd2371447, 25'd3880550, -25'd107793, -25'd1293517, 25'd1149793, 25'd3664964, 25'd3449378}, '{25'd179655, 25'd2479241, 25'd4347654, -25'd35931, 25'd3054137, 25'd287448, 25'd431172, 25'd3125999, -25'd2730758}, '{25'd2443309, 25'd2982275, 25'd4024274, -25'd1113862, -25'd934207, 25'd3593102, -25'd1149793, 25'd2371447, 25'd431172}, '{25'd2982275, 25'd395241, 25'd3449378, -25'd1437241, -25'd1185724, -25'd2119930, -25'd1868413, -25'd1796551, -25'd2694827}, '{25'd4096137, 25'd1365379, 25'd646758, 25'd2443309, 25'd359310, 25'd3054137, 25'd934207, 25'd2658896, -25'd2335516}, '{25'd574896, -25'd3090068, 25'd3125999, -25'd682689, -25'd2335516, 25'd2155861, 25'd4347654, -25'd1976206, -25'd1293517}, '{-25'd862345, -25'd3090068, 25'd1293517, -25'd3197861, -25'd3952412, -25'd970138, 25'd2658896, -25'd431172, -25'd2407378}}, '{'{25'd1904344, 25'd538965, 25'd3161930, 25'd4239861, -25'd3125999, 25'd4060205, 25'd970138, -25'd2407378, -25'd1724689}, '{-25'd2191792, 25'd3557171, 25'd3880550, -25'd3161930, 25'd3161930, -25'd1760620, -25'd3736826, -25'd646758, 25'd574896}, '{-25'd1652827, -25'd1652827, -25'd2982275, -25'd574896, 25'd4096137, 25'd2946344, 25'd3449378, 25'd467103, -25'd3197861}, '{25'd4239861, -25'd3844619, 25'd3593102, 25'd4060205, -25'd2730758, 25'd3377516, 25'd1688758, -25'd646758, 25'd934207}, '{25'd287448, 25'd1832482, 25'd1113862, 25'd718620, -25'd790482, -25'd1329448, -25'd2658896, -25'd179655, -25'd3629033}, '{-25'd2012137, -25'd3341585, -25'd1401310, -25'd359310, -25'd2694827, -25'd898276, -25'd2551103, -25'd2730758, -25'd2048068}, '{25'd2730758, 25'd3557171, 25'd646758, 25'd3772757, -25'd3233792, 25'd2335516, -25'd359310, 25'd1257586, -25'd3557171}, '{25'd1437241, 25'd3090068, -25'd71862, -25'd3054137, -25'd2515172, 25'd898276, 25'd4563240, -25'd1509103, 25'd1293517}, '{-25'd610827, -25'd2299585, 25'd1329448, -25'd2694827, -25'd359310, 25'd2587034, 25'd538965, -25'd1221655, -25'd826414}}, '{'{-25'd1904344, 25'd2515172, -25'd4132068, -25'd1545034, 25'd0, -25'd1760620, -25'd2335516, -25'd2515172, 25'd3161930}, '{25'd4060205, 25'd682689, -25'd898276, 25'd287448, -25'd826414, -25'd3808688, 25'd71862, -25'd3844619, 25'd2694827}, '{25'd2766689, 25'd3161930, -25'd2227723, -25'd682689, 25'd3772757, 25'd1832482, 25'd682689, -25'd1868413, 25'd610827}, '{-25'd3880550, 25'd2802620, -25'd2479241, 25'd3557171, -25'd2119930, 25'd3557171, -25'd1976206, 25'd3341585, 25'd4060205}, '{-25'd1149793, -25'd2407378, -25'd71862, -25'd1329448, -25'd503034, -25'd1760620, -25'd1221655, 25'd1257586, -25'd2694827}, '{25'd610827, 25'd1652827, -25'd4275792, 25'd2910413, 25'd107793, -25'd1580965, 25'd3341585, -25'd3090068, -25'd1473172}, '{25'd2191792, -25'd1688758, -25'd1832482, -25'd1976206, -25'd2479241, 25'd3988343, -25'd3305654, -25'd1976206, 25'd3449378}, '{25'd1293517, 25'd4311723, -25'd1796551, 25'd4275792, -25'd1724689, 25'd3161930, -25'd2155861, -25'd574896, -25'd538965}, '{-25'd4167999, 25'd179655, -25'd1042000, -25'd754551, -25'd1042000, -25'd3700895, -25'd1329448, 25'd4563240, -25'd2838551}}},
    '{'{'{25'd1677203, -25'd3354406, -25'd4269244, 25'd4002416, -25'd3354406, -25'd3278169, -25'd1829676, -25'd2782632, 25'd3735588}, '{25'd2515804, -25'd762365, -25'd3735588, 25'd1448493, 25'd2706396, 25'd800483, 25'd2020267, 25'd1944031, -25'd724247}, '{-25'd4726663, -25'd2363331, -25'd4688544, 25'd952956, 25'd381182, 25'd1181666, -25'd1677203, -25'd2134622, -25'd190591}, '{25'd2515804, 25'd3316287, 25'd2172740, 25'd2592041, -25'd3049460, -25'd2439568, -25'd2592041, -25'd1753439, -25'd2515804}, '{-25'd4879136, -25'd266828, -25'd4383598, 25'd2363331, 25'd1257902, 25'd3049460, 25'd2363331, -25'd2134622, -25'd2896987}, '{25'd3278169, -25'd4421717, 25'd1372257, 25'd419301, 25'd457419, -25'd228709, 25'd343064, 25'd724247, -25'd2210858}, '{25'd2973223, 25'd1410375, -25'd1296020, -25'd4116771, 25'd4040534, -25'd533655, -25'd190591, 25'd800483, -25'd762365}, '{25'd3392524, -25'd3926179, -25'd3849943, 25'd4231125, 25'd3240051, -25'd2020267, -25'd762365, -25'd3506879, 25'd1448493}, '{25'd724247, -25'd2439568, -25'd724247, 25'd2706396, -25'd800483, -25'd2134622, -25'd648010, 25'd2248977, 25'd3735588}}, '{'{-25'd457419, -25'd4879136, 25'd1410375, -25'd2935105, -25'd800483, 25'd648010, -25'd3278169, 25'd3659352, -25'd1143547}, '{25'd952956, -25'd76236, -25'd2935105, -25'd1905912, -25'd3621233, 25'd3392524, 25'd1600966, -25'd3697470, -25'd2439568}, '{-25'd1639085, -25'd2134622, -25'd4459835, 25'd2935105, -25'd3278169, -25'd381182, 25'd3888061, -25'd1905912, 25'd3468760}, '{25'd2782632, 25'd2363331, -25'd4269244, 25'd2515804, 25'd2668277, -25'd4383598, 25'd2363331, -25'd38118, -25'd3735588}, '{25'd3316287, 25'd3087578, 25'd2325213, -25'd1829676, -25'd838601, 25'd3544997, -25'd2973223, -25'd2858869, -25'd724247}, '{-25'd4421717, 25'd2058385, 25'd1524730, -25'd2553923, 25'd2973223, 25'd2592041, 25'd0, -25'd2325213, 25'd2401450}, '{-25'd4612308, -25'd1219784, -25'd4078652, 25'd190591, 25'd381182, 25'd2744514, 25'd2363331, -25'd571774, -25'd2630159}, '{-25'd419301, -25'd2668277, -25'd876720, 25'd2630159, -25'd3964298, -25'd2020267, 25'd3316287, 25'd3087578, -25'd724247}, '{-25'd2706396, -25'd4574190, -25'd3888061, -25'd914838, -25'd266828, -25'd3888061, 25'd2553923, -25'd3735588, -25'd3011342}}, '{'{25'd190591, 25'd3201933, -25'd4116771, 25'd1944031, 25'd3240051, -25'd1982149, -25'd1867794, -25'd800483, 25'd1143547}, '{-25'd4193007, -25'd76236, 25'd495537, 25'd3240051, 25'd3697470, -25'd876720, 25'd2553923, -25'd1486612, -25'd1181666}, '{-25'd571774, 25'd2553923, 25'd762365, -25'd4193007, 25'd1524730, -25'd2058385, 25'd1639085, 25'd2401450, 25'd4040534}, '{-25'd648010, -25'd38118, -25'd991074, 25'd0, -25'd419301, 25'd304946, 25'd648010, 25'd4269244, 25'd2248977}, '{-25'd381182, 25'd3735588, 25'd1753439, -25'd1105429, 25'd800483, -25'd3240051, -25'd3735588, 25'd533655, 25'd3735588}, '{-25'd762365, -25'd4307362, 25'd381182, 25'd2592041, 25'd2401450, -25'd533655, -25'd3125696, -25'd3011342, 25'd1982149}, '{-25'd1448493, -25'd304946, 25'd1448493, 25'd914838, -25'd2592041, 25'd3583115, 25'd3621233, -25'd3278169, 25'd686128}, '{25'd1296020, -25'd343064, -25'd3544997, 25'd1219784, -25'd3240051, -25'd3735588, 25'd3926179, -25'd228709, 25'd1334139}, '{-25'd609892, -25'd1944031, 25'd4002416, 25'd1181666, 25'd2401450, 25'd4383598, 25'd2325213, 25'd533655, 25'd1715321}}},
    '{'{'{-25'd1832092, -25'd1655929, 25'd3347091, 25'd2043487, -25'd2748138, 25'd739883, 25'd458023, 25'd3593719, -25'd2501510}, '{-25'd3488021, 25'd1092209, 25'd2501510, 25'd352325, -25'd2078720, 25'd2712905, 25'd2325347, 25'd563721, -25'd3769881}, '{-25'd1127441, 25'd1444534, -25'd3170928, -25'd1479766, -25'd2677673, -25'd2466277, -25'd810348, 25'd1691162, 25'd634186}, '{-25'd1902557, -25'd2254882, 25'd2431045, 25'd2642440, -25'd1268371, -25'd634186, -25'd3347091, 25'd2360580, 25'd1796859}, '{25'd1832092, -25'd3558486, 25'd3628951, -25'd4086974, 25'd739883, 25'd3065230, 25'd3452788, -25'd4157439, -25'd2748138}, '{-25'd211395, -25'd1655929, -25'd1620697, 25'd3065230, 25'd2431045, -25'd1479766, 25'd3734649, 25'd3910811, 25'd951278}, '{25'd2466277, -25'd4333602, -25'd1902557, -25'd2607208, -25'd1127441, 25'd2078720, 25'd1691162, -25'd3029998, 25'd916046}, '{25'd2959533, -25'd2184417, 25'd2536742, -25'd2466277, 25'd1092209, -25'd2078720, 25'd70465, -25'd4086974, -25'd493255}, '{-25'd2008254, -25'd2607208, 25'd3170928, 25'd2818603, 25'd176163, -25'd2219650, -25'd845581, -25'd3875579, 25'd2008254}}, '{'{25'd4051741, -25'd598953, -25'd2712905, 25'd1655929, -25'd634186, 25'd3981276, 25'd3382323, -25'd563721, 25'd2818603}, '{-25'd2501510, 25'd3523253, -25'd3664184, 25'd2571975, 25'd1444534, -25'd176163, 25'd2818603, -25'd3910811, -25'd2853835}, '{25'd1691162, -25'd2924300, 25'd2043487, -25'd1479766, 25'd3981276, 25'd845581, 25'd704651, -25'd880813, 25'd880813}, '{25'd1832092, -25'd352325, -25'd1937789, 25'd2078720, 25'd634186, 25'd1409301, 25'd2254882, -25'd598953, 25'd3734649}, '{-25'd739883, -25'd4227904, 25'd2994765, 25'd493255, 25'd1514999, 25'd951278, 25'd3488021, -25'd775116, 25'd3065230}, '{-25'd3805114, -25'd2325347, 25'd1409301, 25'd0, -25'd1409301, 25'd3558486, 25'd3347091, -25'd1902557, -25'd3029998}, '{25'd3840346, -25'd3840346, 25'd704651, -25'd2431045, -25'd35233, 25'd1162674, -25'd1902557, -25'd3452788, 25'd2466277}, '{25'd0, -25'd2712905, 25'd2149185, 25'd739883, 25'd387558, -25'd35233, 25'd2431045, -25'd2677673, 25'd1374069}, '{25'd3628951, 25'd35233, -25'd1021743, 25'd1303604, -25'd3382323, 25'd1479766, 25'd1197906, -25'd1655929, -25'd1973022}}, '{'{-25'd35233, -25'd2008254, 25'd1479766, -25'd986511, 25'd1374069, -25'd3805114, -25'd2571975, 25'd458023, 25'd2571975}, '{25'd1761627, -25'd2818603, 25'd1374069, 25'd1691162, 25'd281860, -25'd1514999, 25'd2818603, 25'd4086974, -25'd4192672}, '{25'd563721, 25'd4474532, 25'd2501510, -25'd3488021, 25'd1056976, 25'd211395, 25'd3981276, 25'd880813, 25'd4051741}, '{-25'd3734649, 25'd1867324, 25'd4474532, 25'd3065230, 25'd2113952, 25'd1796859, -25'd3241393, -25'd2113952, -25'd2783370}, '{-25'd3699416, -25'd2501510, -25'd1761627, 25'd2818603, -25'd458023, -25'd1021743, 25'd1585464, 25'd2853835, 25'd3311858}, '{25'd3311858, -25'd3769881, -25'd3311858, -25'd775116, -25'd3523253, 25'd140930, 25'd2466277, -25'd986511, -25'd3382323}, '{-25'd1585464, -25'd634186, -25'd1550232, -25'd1092209, 25'd1902557, 25'd2889068, -25'd669418, 25'd1092209, 25'd211395}, '{25'd2431045, 25'd2818603, 25'd3628951, -25'd3910811, -25'd3628951, 25'd4227904, 25'd3135696, 25'd2818603, 25'd845581}, '{25'd3910811, 25'd2078720, 25'd3769881, 25'd3311858, -25'd1585464, 25'd3135696, 25'd4227904, -25'd3311858, -25'd986511}}},
    '{'{'{-25'd1099603, 25'd1620468, -25'd1620468, -25'd1504720, -25'd57874, -25'd983856, -25'd3530306, 25'd231495, -25'd3472432}, '{-25'd5035026, -25'd2546450, 25'd2372828, -25'd5555891, -25'd2720072, -25'd4687783, -25'd5208648, -25'd6018882, -25'd3761801}, '{-25'd5382269, -25'd4803531, -25'd4803531, -25'd4282666, 25'd3646053, 25'd4166918, 25'd2372828, 25'd983856, 25'd1620468}, '{-25'd231495, -25'd3819675, 25'd2604324, 25'd4340540, -25'd694486, -25'd1215351, 25'd5150774, 25'd3646053, -25'd636612}, '{25'd1504720, -25'd173622, -25'd578739, -25'd1388973, 25'd6134629, 25'd5555891, 25'd2835819, 25'd4456287, 25'd1099603}, '{25'd3009441, 25'd5150774, 25'd2257081, 25'd4166918, -25'd173622, 25'd3819675, 25'd868108, -25'd1736216, 25'd2372828}, '{25'd1909837, 25'd520865, -25'd2199207, 25'd347243, 25'd3414558, 25'd4109044, 25'd4572035, 25'd1331099, -25'd3067315}, '{-25'd2257081, 25'd1851964, 25'd4977152, -25'd1620468, 25'd2488576, -25'd405117, 25'd4456287, 25'd2141333, 25'd3414558}, '{25'd3125189, 25'd5150774, 25'd925982, -25'd1851964, -25'd983856, -25'd2083459, 25'd5440143, -25'd2662198, -25'd173622}}, '{'{-25'd3877549, -25'd2083459, -25'd6134629, 25'd2546450, 25'd2141333, 25'd3009441, -25'd1273225, 25'd925982, 25'd1388973}, '{25'd925982, -25'd2314955, -25'd5671639, 25'd578739, -25'd2141333, -25'd4687783, -25'd3993297, -25'd4340540, -25'd4919278}, '{25'd1504720, -25'd1099603, -25'd3588179, -25'd694486, 25'd173622, -25'd4109044, -25'd1794090, -25'd3472432, 25'd2430702}, '{25'd3125189, 25'd752360, 25'd0, -25'd173622, 25'd694486, -25'd2141333, 25'd405117, 25'd4456287, -25'd1678342}, '{-25'd2314955, 25'd1678342, -25'd752360, -25'd1099603, 25'd7349981, 25'd7002737, 25'd4514161, -25'd1794090, 25'd3819675}, '{-25'd2662198, 25'd3761801, 25'd578739, 25'd5382269, 25'd2199207, 25'd289369, 25'd462991, 25'd868108, 25'd4803531}, '{25'd1851964, -25'd2546450, -25'd1388973, 25'd2720072, 25'd2314955, 25'd3819675, 25'd5613765, -25'd1909837, 25'd4745657}, '{-25'd1099603, 25'd2314955, 25'd810234, 25'd1041730, -25'd1273225, -25'd2372828, 25'd4745657, 25'd3067315, 25'd4629909}, '{25'd578739, -25'd925982, 25'd4861404, -25'd1678342, 25'd4340540, -25'd1504720, 25'd5671639, -25'd2083459, -25'd2083459}}, '{'{-25'd1388973, 25'd1851964, -25'd4282666, -25'd4109044, 25'd173622, -25'd3935423, -25'd5555891, 25'd2199207, 25'd1620468}, '{-25'd5440143, -25'd3125189, 25'd289369, -25'd4166918, -25'd3819675, -25'd4398414, -25'd694486, -25'd2777945, -25'd1446847}, '{-25'd4282666, -25'd3819675, -25'd1967711, 25'd1041730, 25'd3530306, -25'd694486, 25'd3298810, -25'd5035026, -25'd2893693}, '{25'd578739, 25'd115748, 25'd925982, -25'd636612, -25'd1794090, 25'd4051170, 25'd173622, -25'd1504720, -25'd4224792}, '{25'd462991, 25'd5035026, 25'd2141333, 25'd231495, -25'd115748, 25'd5498017, -25'd2083459, 25'd2257081, 25'd3125189}, '{-25'd2430702, 25'd694486, 25'd4919278, -25'd462991, 25'd6655494, 25'd4166918, 25'd347243, 25'd1273225, 25'd1099603}, '{25'd4051170, 25'd1678342, 25'd5208648, -25'd1736216, 25'd4572035, 25'd5729512, 25'd3935423, -25'd173622, -25'd2314955}, '{-25'd868108, -25'd1215351, 25'd2314955, 25'd4861404, 25'd5208648, 25'd4109044, 25'd1736216, -25'd3240936, -25'd1215351}, '{25'd1099603, 25'd1157477, 25'd694486, 25'd2430702, -25'd57874, -25'd289369, 25'd1620468, -25'd810234, -25'd2546450}}},
    '{'{'{-25'd1680677, 25'd3738648, -25'd1612078, 25'd3738648, -25'd926087, -25'd3567150, 25'd1406280, 25'd1474879, 25'd4321740}, '{25'd34300, -25'd3189856, 25'd1920773, 25'd3944445, -25'd720290, -25'd3738648, 25'd3807247, 25'd3395653, -25'd2092271}, '{25'd4150242, -25'd2881160, -25'd3738648, 25'd2229469, -25'd3807247, 25'd3841546, -25'd2469566, 25'd1166184, -25'd1955073}, '{25'd3361353, 25'd1989372, 25'd1131884, 25'd4150242, 25'd137198, 25'd3121257, -25'd2092271, -25'd2984058, -25'd1749276}, '{25'd651691, -25'd2160870, 25'd1680677, 25'd34300, 25'd2435266, 25'd4218841, 25'd857488, -25'd583092, -25'd1269082}, '{-25'd926087, -25'd1955073, -25'd2092271, 25'd994686, 25'd3086957, 25'd4253141, 25'd4356039, 25'd823189, -25'd2057971}, '{25'd2435266, -25'd3738648, -25'd3361353, -25'd2709662, 25'd1440580, 25'd857488, 25'd137198, -25'd342995, -25'd4218841}, '{-25'd3567150, 25'd1680677, -25'd823189, -25'd994686, 25'd3841546, -25'd3052657, -25'd1097585, -25'd2778261, -25'd3292754}, '{-25'd68599, 25'd3567150, -25'd2469566, -25'd754589, 25'd2263768, 25'd205797, 25'd411594, 25'd1852174, -25'd651691}}, '{'{25'd2469566, -25'd2160870, 25'd2229469, -25'd685990, 25'd3635749, 25'd891788, -25'd1371981, 25'd3018358, -25'd171498}, '{-25'd1612078, -25'd3978745, 25'd1063285, -25'd1509179, 25'd3464252, -25'd2812561, 25'd3292754, -25'd2881160, 25'd3292754}, '{25'd4321740, 25'd1577778, -25'd3807247, 25'd3292754, -25'd2572464, -25'd342995, -25'd4081643, 25'd274396, 25'd2195169}, '{25'd3464252, 25'd377295, 25'd4047344, -25'd2984058, -25'd2572464, -25'd3910146, -25'd3498551, -25'd2126570, -25'd3121257}, '{25'd1543479, 25'd1680677, -25'd445894, -25'd3807247, -25'd651691, 25'd2641063, 25'd1234783, 25'd411594, 25'd4321740}, '{25'd2023672, -25'd1509179, 25'd720290, 25'd685990, -25'd3155556, 25'd1131884, 25'd2984058, -25'd274396, 25'd4218841}, '{25'd2366667, 25'd2160870, -25'd411594, -25'd3086957, 25'd2675363, 25'd2400967, -25'd788889, -25'd3532851, 25'd583092}, '{-25'd3189856, 25'd4321740, 25'd4150242, 25'd823189, 25'd3189856, -25'd685990, 25'd1337681, 25'd788889, 25'd3910146}, '{-25'd754589, -25'd3498551, -25'd308696, -25'd1680677, -25'd891788, 25'd960387, -25'd137198, -25'd2160870, 25'd3841546}}, '{'{25'd4081643, -25'd823189, 25'd1749276, 25'd377295, 25'd3601450, -25'd1166184, 25'd3635749, -25'd788889, -25'd2023672}, '{25'd3910146, 25'd3327054, -25'd4115943, -25'd960387, 25'd1474879, 25'd1371981, -25'd685990, -25'd102899, 25'd926087}, '{-25'd1371981, 25'd3841546, -25'd3361353, -25'd3121257, -25'd3189856, 25'd3738648, -25'd2984058, 25'd1783575, 25'd1783575}, '{-25'd3429952, 25'd2435266, 25'd2229469, -25'd1749276, 25'd308696, -25'd685990, 25'd2195169, -25'd926087, 25'd514493}, '{25'd2915459, -25'd583092, -25'd2984058, 25'd514493, 25'd891788, -25'd2366667, 25'd4321740, 25'd2195169, 25'd2709662}, '{25'd548792, 25'd1543479, -25'd3498551, -25'd514493, 25'd4047344, -25'd3155556, -25'd994686, 25'd3601450, 25'd68599}, '{25'd3429952, 25'd2915459, -25'd4047344, -25'd617391, -25'd3018358, -25'd2023672, -25'd2881160, 25'd2915459, 25'd0}, '{-25'd3841546, 25'd4047344, -25'd3327054, -25'd514493, -25'd960387, 25'd651691, 25'd2092271, 25'd3772947, 25'd1097585}, '{25'd514493, 25'd1303382, -25'd4287440, 25'd3978745, -25'd2092271, -25'd3052657, 25'd4115943, 25'd102899, 25'd3052657}}},
    '{'{'{-25'd3150513, -25'd2737946, -25'd1650269, 25'd150024, -25'd1125183, 25'd1537750, 25'd3563080, 25'd2175354, -25'd862640}, '{25'd2587921, -25'd2587921, 25'd4763276, 25'd2325379, 25'd1462738, -25'd1462738, 25'd1687775, -25'd637604, 25'd4388215}, '{25'd1762787, 25'd150024, 25'd2175354, 25'd1500244, 25'd4725770, -25'd75012, 25'd712616, 25'd1800293, 25'd3188019}, '{-25'd1312714, -25'd1125183, 25'd675110, 25'd3825623, 25'd4163178, 25'd3300538, -25'd787628, -25'd3900635, 25'd1500244}, '{25'd487579, 25'd4313202, -25'd3675599, 25'd112518, 25'd1987824, 25'd2362885, 25'd4763276, -25'd337555, -25'd2025330}, '{25'd2700440, -25'd2737946, -25'd3188019, 25'd4050660, 25'd3675599, -25'd1687775, 25'd3413056, 25'd3600586, 25'd1725281}, '{25'd1650269, 25'd4125672, 25'd4463227, -25'd75012, 25'd1125183, -25'd712616, -25'd1537750, 25'd3938141, 25'd225037}, '{25'd112518, -25'd3150513, 25'd3938141, 25'd2100342, -25'd1425232, 25'd2400391, -25'd2625428, -25'd75012, 25'd2662934}, '{-25'd712616, -25'd787628, 25'd787628, 25'd2550415, -25'd1125183, 25'd4313202, -25'd1462738, -25'd1762787, -25'd1800293}}, '{'{-25'd2512909, 25'd1387726, -25'd1237702, -25'd2400391, -25'd2175354, -25'd2362885, 25'd3675599, -25'd3600586, 25'd1200195}, '{-25'd3863129, 25'd1087677, 25'd3300538, -25'd1162689, 25'd375061, 25'd187531, 25'd2437897, 25'd3375550, -25'd3825623}, '{-25'd1612763, -25'd3713105, -25'd2737946, 25'd3863129, -25'd1762787, 25'd2400391, 25'd4463227, 25'd375061, 25'd637604}, '{25'd4425721, -25'd150024, -25'd300049, -25'd1575257, -25'd1200195, -25'd3563080, 25'd300049, -25'd2287873, 25'd412567}, '{-25'd300049, -25'd337555, -25'd2362885, -25'd2475403, 25'd4425721, -25'd3525574, 25'd4425721, 25'd3750611, 25'd1125183}, '{25'd3863129, -25'd1162689, -25'd1987824, -25'd3900635, 25'd4200684, 25'd1987824, 25'd4613251, 25'd2437897, -25'd1687775}, '{25'd3037995, -25'd3000489, -25'd862640, -25'd3037995, 25'd2625428, -25'd900147, 25'd3225525, -25'd2662934, -25'd900147}, '{25'd2587921, -25'd2175354, -25'd3600586, -25'd2175354, 25'd1875305, 25'd1012665, -25'd75012, 25'd1912812, 25'd1762787}, '{-25'd2925476, -25'd2362885, -25'd2587921, 25'd2475403, 25'd4050660, 25'd1237702, 25'd862640, 25'd412567, 25'd225037}}, '{'{-25'd3225525, 25'd2700440, 25'd1800293, -25'd1837799, -25'd1800293, -25'd2062836, -25'd3675599, 25'd2025330, 25'd0}, '{-25'd2587921, 25'd1012665, -25'd112518, 25'd3413056, 25'd1500244, -25'd2362885, -25'd675110, -25'd3375550, -25'd787628}, '{25'd1875305, -25'd1950318, -25'd2175354, -25'd900147, 25'd450073, -25'd562592, 25'd1462738, 25'd4350709, 25'd2400391}, '{-25'd825134, 25'd4613251, 25'd2100342, -25'd2325379, 25'd4313202, -25'd1537750, -25'd1650269, -25'd2737946, -25'd525086}, '{-25'd1537750, 25'd4163178, -25'd1162689, -25'd2025330, -25'd2100342, 25'd3037995, 25'd2250367, -25'd1875305, 25'd4463227}, '{25'd1950318, 25'd675110, 25'd4013154, 25'd975159, 25'd0, 25'd1162689, 25'd4388215, -25'd1012665, -25'd1275208}, '{-25'd3863129, -25'd1875305, 25'd825134, -25'd1125183, 25'd3113007, 25'd4125672, 25'd1650269, -25'd3188019, 25'd4388215}, '{-25'd1612763, 25'd2212860, 25'd4575745, 25'd1162689, 25'd2287873, -25'd637604, -25'd3413056, -25'd1987824, 25'd300049}, '{25'd2550415, -25'd1725281, -25'd112518, 25'd4088166, 25'd4763276, -25'd3750611, -25'd1462738, 25'd1800293, 25'd4125672}}},
    '{'{'{25'd925283, -25'd3772308, -25'd1281161, 25'd3060551, 25'd35588, 25'd3096139, -25'd177939, -25'd3629956, -25'd2384383}, '{-25'd1565864, 25'd3736720, -25'd3416430, 25'd2740261, -25'd1281161, -25'd2811437, 25'd4270537, 25'd604993, 25'd2206444}, '{-25'd1067634, -25'd3914659, 25'd4021422, 25'd533817, 25'd2491147, -25'd2491147, 25'd4270537, 25'd1850566, 25'd177939}, '{25'd2384383, 25'd3985834, 25'd889695, 25'd1637039, 25'd1743803, -25'd4021422, -25'd569405, 25'd1209985, 25'd3914659}, '{25'd1957329, 25'd711756, 25'd3274078, -25'd284702, 25'd3452017, -25'd2064093, -25'd3060551, -25'd4092598, 25'd1459100}, '{-25'd3665544, -25'd1423512, -25'd2526734, -25'd1494688, -25'd1352337, 25'd1352337, 25'd1743803, 25'd818520, -25'd1814978}, '{-25'd2313207, -25'd1423512, -25'd960871, 25'd3701132, -25'd4234949, 25'd1281161, -25'd3772308, 25'd3096139, -25'd2028505}, '{-25'd4377300, 25'd3309666, 25'd996459, 25'd1601451, 25'd782932, 25'd355878, 25'd355878, 25'd854107, 25'd2206444}, '{25'd996459, 25'd2313207, 25'd3736720, -25'd4128186, 25'd676168, 25'd925283, -25'd533817, 25'd3416430, 25'd3950247}}, '{'{25'd1601451, -25'd2847025, 25'd747344, 25'd1672627, 25'd1921742, 25'd3843483, -25'd2313207, 25'd676168, 25'd1850566}, '{-25'd2348795, 25'd2882612, 25'd2918200, 25'd2526734, -25'd2847025, -25'd142351, -25'd1779390, 25'd2953788, -25'd1459100}, '{25'd498229, -25'd3345254, 25'd1352337, 25'd3843483, -25'd2384383, 25'd2313207, 25'd320290, 25'd1601451, -25'd3060551}, '{-25'd142351, -25'd355878, -25'd284702, 25'd996459, -25'd2953788, -25'd3309666, -25'd1530276, -25'd2704673, -25'd1352337}, '{-25'd1103222, 25'd2989376, -25'd1672627, 25'd320290, 25'd1387924, -25'd2242032, 25'd2953788, 25'd640581, -25'd1708215}, '{25'd142351, -25'd1637039, 25'd3558781, -25'd3879071, 25'd2669086, -25'd2704673, -25'd2918200, -25'd960871, 25'd71176}, '{25'd3807895, -25'd676168, -25'd960871, -25'd2170856, -25'd533817, -25'd249115, 25'd1174398, 25'd2597910, -25'd1032046}, '{25'd4057010, 25'd4163773, -25'd3950247, 25'd3879071, 25'd1601451, 25'd4341713, 25'd2989376, 25'd1423512, 25'd3843483}, '{25'd676168, 25'd3452017, 25'd2847025, 25'd996459, 25'd3274078, 25'd4199361, -25'd3380842, 25'd3060551, 25'd3060551}}, '{'{25'd2277620, 25'd427054, 25'd1494688, -25'd2384383, 25'd1957329, 25'd4021422, -25'd3558781, -25'd3380842, 25'd1209985}, '{-25'd3096139, -25'd2384383, -25'd3345254, 25'd1992917, 25'd854107, 25'd2597910, 25'd996459, 25'd1494688, -25'd2099681}, '{25'd2775849, -25'd854107, 25'd3487605, -25'd4057010, 25'd213527, 25'd106763, 25'd3629956, -25'd2099681, -25'd2562322}, '{-25'd2277620, -25'd106763, -25'd747344, -25'd3416430, -25'd4555239, 25'd2028505, -25'd3345254, 25'd2597910, 25'd3914659}, '{25'd1957329, 25'd2669086, -25'd3131727, 25'd1565864, -25'd1886154, 25'd3202903, -25'd604993, -25'd1921742, -25'd2348795}, '{25'd2170856, 25'd2455559, 25'd3950247, -25'd1067634, 25'd3452017, -25'd3024964, 25'd569405, 25'd391466, -25'd3807895}, '{25'd854107, 25'd3309666, 25'd391466, -25'd569405, -25'd4377300, -25'd2740261, -25'd1032046, -25'd320290, -25'd2526734}, '{-25'd177939, 25'd1601451, 25'd249115, -25'd3238490, 25'd1032046, -25'd1565864, -25'd604993, 25'd2847025, 25'd3701132}, '{-25'd142351, -25'd3950247, -25'd2633498, 25'd3060551, 25'd1387924, -25'd462641, 25'd3558781, -25'd4128186, 25'd1494688}}},
    '{'{'{25'd3925776, 25'd4000553, -25'd3065844, 25'd598214, 25'd822544, -25'd3477116, 25'd2018971, -25'd2131136, -25'd672990}, '{-25'd897320, 25'd2729349, -25'd224330, -25'd1757252, 25'd486048, -25'd3664058, -25'd1196427, 25'd1981582, 25'd1682476}, '{25'd3888388, 25'd3140621, -25'd710379, 25'd1607699, 25'd1794641, 25'd3252786, -25'd1794641, 25'd2131136, 25'd261718}, '{25'd897320, 25'd4112718, 25'd3514505, -25'd2542408, 25'd1383369, 25'd1383369, 25'd2729349, -25'd3215398, -25'd2916291}, '{-25'd2505019, 25'd411272, -25'd822544, -25'd1682476, 25'd4037941, -25'd1757252, -25'd2467631, 25'd672990, 25'd3402339}, '{25'd2243301, 25'd1719864, -25'd3215398, 25'd186942, 25'd785155, 25'd3215398, 25'd1345980, 25'd3925776, -25'd112165}, '{25'd2617184, -25'd1420757, -25'd3065844, 25'd2205912, 25'd3364951, 25'd710379, 25'd373883, 25'd1719864, -25'd1009485}, '{25'd3402339, 25'd934709, 25'd3551893, 25'd4187495, -25'd1009485, -25'd37388, -25'd1009485, -25'd3589281, 25'd1009485}, '{-25'd1383369, 25'd3028456, -25'd1271204, -25'd822544, -25'd2878903, -25'd448660, -25'd3925776, -25'd1869417, -25'd1719864}}, '{'{-25'd2243301, 25'd635602, -25'd2654573, -25'd3589281, 25'd1009485, 25'd186942, -25'd3439728, 25'd3028456, -25'd785155}, '{-25'd3290174, -25'd3963165, -25'd1869417, -25'd1832029, 25'd3402339, -25'd2654573, -25'd3290174, -25'd2205912, -25'd4710932}, '{25'd2355466, -25'd1084262, 25'd1345980, -25'd2056359, -25'd3364951, 25'd3215398, 25'd747767, 25'd411272, 25'd1159039}, '{-25'd224330, -25'd4150106, -25'd3252786, -25'd4785708, 25'd897320, 25'd1495534, 25'd1009485, -25'd1944194, 25'd3551893}, '{25'd3589281, 25'd1832029, 25'd149553, -25'd2766738, -25'd4449213, -25'd4411825, 25'd2093747, -25'd1645087, 25'd2766738}, '{-25'd4486602, 25'd2318077, -25'd3065844, -25'd3551893, -25'd2916291, -25'd4000553, -25'd2654573, 25'd635602, 25'd2392854}, '{25'd224330, -25'd2131136, -25'd1046874, 25'd1009485, -25'd3327563, -25'd112165, 25'd224330, -25'd3178009, -25'd1383369}, '{25'd1009485, 25'd37388, -25'd4224883, -25'd1757252, 25'd4000553, 25'd747767, 25'd2729349, -25'd2505019, 25'd1196427}, '{25'd1682476, -25'd1645087, 25'd2355466, 25'd1645087, 25'd2355466, -25'd2355466, -25'd1196427, 25'd1607699, -25'd1832029}}, '{'{-25'd1906806, 25'd710379, -25'd1682476, 25'd2804126, -25'd3215398, -25'd336495, 25'd1196427, -25'd2841514, -25'd3103233}, '{-25'd635602, -25'd373883, -25'd4187495, 25'd1084262, -25'd4187495, -25'd3215398, 25'd2766738, -25'd859932, 25'd1607699}, '{25'd112165, 25'd74777, -25'd2467631, -25'd747767, 25'd186942, -25'd523437, -25'd3963165, 25'd2318077, -25'd560825}, '{25'd3439728, 25'd1757252, -25'd4000553, -25'd897320, -25'd3963165, -25'd859932, -25'd2280689, 25'd2916291, -25'd3252786}, '{25'd411272, -25'd3551893, -25'd1383369, 25'd3813611, -25'd897320, -25'd2243301, 25'd3477116, 25'd2093747, -25'd2804126}, '{-25'd1570311, 25'd2131136, -25'd2916291, -25'd2018971, -25'd2654573, -25'd2355466, -25'd4598767, -25'd2392854, -25'd4411825}, '{25'd4411825, 25'd3738835, -25'd299107, -25'd2392854, -25'd1944194, 25'd3551893, -25'd261718, -25'd373883, -25'd2841514}, '{25'd3477116, 25'd1159039, -25'd1682476, -25'd1869417, -25'd3215398, -25'd1981582, 25'd934709, -25'd3664058, 25'd672990}, '{25'd747767, 25'd2505019, 25'd2168524, -25'd3813611, -25'd1495534, 25'd3776223, -25'd2991068, 25'd3065844, 25'd336495}}},
    '{'{'{-25'd845693, 25'd1434002, -25'd1323694, -25'd404462, -25'd1801694, -25'd3419542, 25'd1139847, -25'd1470771, -25'd3713697}, '{25'd2684157, -25'd3713697, -25'd3088619, 25'd4154928, 25'd3125388, 25'd3713697, 25'd3971082, -25'd2169387, 25'd2022310}, '{-25'd4302005, 25'd2647388, -25'd992770, -25'd3309235, 25'd992770, -25'd4302005, -25'd3382773, 25'd1801694, 25'd3493081}, '{-25'd404462, 25'd2684157, -25'd36769, -25'd882463, 25'd2941542, 25'd1617848, 25'd2059079, -25'd3934312, 25'd3676927}, '{25'd1654617, -25'd1691387, -25'd367693, -25'd1581079, 25'd3419542, -25'd1581079, 25'd1434002, 25'd845693, -25'd661847}, '{25'd1139847, 25'd2132618, 25'd1360463, -25'd3860774, -25'd2794465, -25'd147077, -25'd3603389, 25'd2757696, 25'd2059079}, '{-25'd294154, -25'd1764925, -25'd1764925, -25'd4485851, 25'd808924, -25'd3272465, 25'd110308, 25'd3787235, -25'd625078}, '{-25'd3419542, -25'd3971082, -25'd3309235, 25'd257385, -25'd2279695, -25'd1764925, -25'd919232, -25'd257385, -25'd3971082}, '{25'd441231, -25'd4191697, -25'd1507540, -25'd441231, -25'd3640158, -25'd441231, -25'd2022310, 25'd147077, -25'd2169387}}, '{'{-25'd551539, 25'd3015080, -25'd1654617, -25'd4596159, 25'd1176617, -25'd73539, 25'd845693, -25'd36769, -25'd3824005}, '{-25'd4706467, -25'd4118159, 25'd3603389, 25'd478001, -25'd404462, 25'd441231, 25'd2022310, 25'd514770, 25'd2941542}, '{-25'd808924, 25'd3824005, -25'd367693, 25'd1654617, -25'd772155, 25'd919232, -25'd220616, -25'd3456312, 25'd1985541}, '{25'd2169387, -25'd1029540, 25'd3456312, 25'd2206156, -25'd1912002, -25'd1875233, -25'd4081389, -25'd3419542, -25'd1617848}, '{25'd1360463, -25'd2022310, 25'd3309235, 25'd698616, -25'd2978311, -25'd330923, -25'd3566620, 25'd367693, -25'd3051850}, '{25'd183846, 25'd257385, 25'd2757696, 25'd3824005, 25'd3897543, -25'd1654617, 25'd147077, -25'd73539, -25'd4596159}, '{25'd3125388, -25'd3309235, 25'd3309235, -25'd330923, -25'd4191697, 25'd3088619, -25'd4412313, -25'd625078, -25'd4706467}, '{-25'd4412313, -25'd1691387, 25'd2132618, 25'd2941542, -25'd2904773, -25'd3676927, -25'd3640158, 25'd992770, -25'd4228467}, '{-25'd3603389, 25'd73539, -25'd1213386, -25'd3676927, -25'd330923, -25'd1029540, 25'd1801694, 25'd2279695, 25'd1286925}}, '{'{25'd2242926, 25'd551539, 25'd1985541, -25'd3125388, 25'd330923, 25'd1139847, -25'd2647388, 25'd3235696, -25'd4338774}, '{-25'd2353234, 25'd3346004, -25'd2353234, -25'd3971082, -25'd36769, 25'd36769, 25'd1139847, 25'd2242926, 25'd1948772}, '{-25'd3272465, 25'd2573849, -25'd110308, -25'd4228467, -25'd1470771, -25'd2132618, 25'd882463, 25'd294154, -25'd2059079}, '{25'd992770, -25'd1139847, 25'd3015080, 25'd2353234, 25'd2831234, 25'd2831234, 25'd110308, -25'd1985541, 25'd3750466}, '{-25'd2757696, 25'd0, 25'd1764925, 25'd3456312, 25'd1176617, 25'd2831234, 25'd625078, 25'd4007851, 25'd698616}, '{-25'd2390003, 25'd2794465, -25'd1948772, -25'd1213386, -25'd220616, 25'd3934312, 25'd1176617, 25'd1764925, 25'd478001}, '{-25'd367693, 25'd3529850, -25'd1397232, 25'd661847, 25'd1948772, -25'd551539, 25'd1176617, 25'd2390003, -25'd110308}, '{-25'd808924, 25'd2169387, -25'd330923, 25'd3198927, 25'd1985541, -25'd4412313, -25'd2426772, -25'd1213386, -25'd2941542}, '{-25'd625078, -25'd4265236, -25'd257385, -25'd625078, 25'd2831234, 25'd1544310, 25'd3529850, -25'd404462, 25'd3382773}}},
    '{'{'{25'd2914792, -25'd705192, 25'd1222332, -25'd423115, 25'd4090111, -25'd94026, -25'd3102843, 25'd141038, -25'd2632715}, '{-25'd752204, 25'd2068562, 25'd188051, -25'd188051, -25'd2632715, 25'd3008817, -25'd3243881, 25'd5077379, -25'd235064}, '{25'd2350639, -25'd2867779, -25'd4231150, -25'd1833498, -25'd893243, -25'd987268, 25'd3196869, 25'd5970622, 25'd2773754}, '{25'd1974536, -25'd2162588, -25'd4043098, -25'd2726741, -25'd4983354, -25'd2726741, 25'd4466213, 25'd5547507, -25'd2021549}, '{25'd3196869, -25'd3761022, 25'd188051, -25'd4466213, -25'd4513226, -25'd1645447, -25'd2444664, 25'd564153, -25'd2303626}, '{25'd3902060, -25'd2444664, 25'd1974536, 25'd3102843, -25'd5171405, -25'd5218418, -25'd2726741, -25'd282077, -25'd2021549}, '{25'd5500494, 25'd1551422, -25'd1034281, -25'd987268, -25'd1457396, -25'd3290894, -25'd3619984, 25'd2397651, -25'd1316358}, '{-25'd517141, -25'd2209600, 25'd329089, 25'd4701277, -25'd564153, 25'd1363370, -25'd846230, 25'd3808035, 25'd5641533}, '{25'd4513226, 25'd611166, -25'd2162588, -25'd517141, 25'd2820766, 25'd4560239, -25'd2491677, 25'd2256613, 25'd3855047}}, '{'{25'd2115575, -25'd423115, -25'd2726741, 25'd1974536, 25'd987268, -25'd1457396, 25'd2444664, -25'd1927524, 25'd235064}, '{25'd1316358, 25'd2726741, -25'd3478945, 25'd3384920, 25'd705192, -25'd2914792, 25'd376102, -25'd329089, 25'd1551422}, '{25'd799217, 25'd3290894, -25'd3666996, 25'd2115575, 25'd1598434, 25'd1927524, 25'd4372188, 25'd987268, 25'd2820766}, '{-25'd2256613, -25'd3290894, -25'd2961805, -25'd4090111, 25'd1222332, 25'd1081294, -25'd987268, -25'd1269345, -25'd752204}, '{25'd4795303, -25'd2632715, -25'd1457396, -25'd2115575, -25'd2726741, -25'd94026, -25'd2303626, -25'd2632715, 25'd3902060}, '{25'd3337907, 25'd1645447, 25'd2115575, -25'd893243, -25'd5124392, -25'd4936341, -25'd3761022, 25'd4607252, 25'd4654265}, '{-25'd1457396, -25'd2115575, 25'd1786485, -25'd4701277, -25'd1175319, -25'd2538690, 25'd3196869, 25'd1739473, -25'd3714009}, '{25'd3949073, -25'd1974536, -25'd658179, -25'd1551422, 25'd376102, 25'd1363370, 25'd1739473, 25'd3243881, -25'd376102}, '{-25'd1316358, 25'd3902060, 25'd3855047, 25'd1974536, -25'd1316358, 25'd2444664, 25'd4043098, 25'd4513226, 25'd1974536}}, '{'{-25'd611166, 25'd3149856, -25'd3949073, -25'd4466213, -25'd1269345, 25'd282077, -25'd470128, 25'd3808035, 25'd3102843}, '{25'd3525958, 25'd3384920, -25'd2397651, -25'd2350639, 25'd705192, -25'd470128, 25'd4278162, 25'd0, 25'd376102}, '{-25'd1974536, -25'd564153, 25'd3478945, -25'd752204, 25'd2914792, 25'd3008817, 25'd4560239, 25'd1410383, 25'd2773754}, '{-25'd3290894, 25'd1363370, -25'd4325175, 25'd3102843, 25'd752204, 25'd1927524, 25'd188051, 25'd4748290, -25'd1034281}, '{-25'd893243, -25'd1222332, 25'd1316358, -25'd1175319, 25'd564153, -25'd329089, -25'd3008817, 25'd329089, 25'd1363370}, '{25'd3761022, -25'd705192, 25'd2303626, 25'd235064, 25'd235064, 25'd1739473, -25'd3384920, -25'd2162588, -25'd329089}, '{-25'd3337907, -25'd47013, 25'd2961805, 25'd611166, -25'd5218418, -25'd3525958, -25'd1645447, -25'd2397651, -25'd2538690}, '{25'd2914792, -25'd752204, -25'd752204, -25'd2867779, -25'd4560239, -25'd3996086, -25'd705192, -25'd329089, -25'd2209600}, '{25'd2491677, 25'd752204, 25'd3149856, 25'd611166, 25'd1504409, -25'd2350639, -25'd1786485, 25'd1786485, -25'd188051}}},
    '{'{'{25'd2463418, -25'd197073, 25'd837562, 25'd2759028, -25'd2709760, 25'd1724393, -25'd640489, -25'd4187811, 25'd4089274}, '{25'd3941469, 25'd1379514, -25'd1182441, -25'd1724393, -25'd886830, 25'd1872198, -25'd2906833, -25'd886830, -25'd689757}, '{-25'd3251712, 25'd2167808, -25'd4040005, 25'd3153175, -25'd2217076, 25'd3547322, -25'd246342, 25'd4384884, -25'd1034636}, '{-25'd2414150, 25'd295610, -25'd2561955, -25'd837562, 25'd3005370, -25'd2217076, 25'd1330246, -25'd3842932, 25'd3941469}, '{25'd4286347, -25'd1625856, -25'd344879, -25'd3251712, -25'd1773661, 25'd886830, 25'd886830, 25'd3941469, 25'd3300980}, '{25'd3744395, -25'd985367, -25'd3695127, 25'd492684, 25'd4138542, 25'd1970734, -25'd4040005, -25'd3990737, -25'd3202443}, '{-25'd1231709, -25'd1133172, -25'd3547322, -25'd2956102, -25'd3744395, 25'd344879, 25'd1625856, -25'd3941469, -25'd3941469}, '{25'd2611223, 25'd1576588, -25'd1625856, -25'd3498054, -25'd1182441, -25'd295610, -25'd3399517, -25'd4532689, 25'd3793664}, '{-25'd2759028, 25'd1231709, -25'd2906833, 25'd1083904, -25'd2906833, -25'd689757, -25'd4089274, -25'd886830, -25'd1724393}}, '{'{-25'd3103907, -25'd1724393, 25'd3448785, 25'd2906833, -25'd2512686, -25'd1970734, 25'd2561955, 25'd1182441, -25'd1182441}, '{-25'd197073, 25'd739025, -25'd3054638, 25'd3498054, 25'd1034636, 25'd1133172, 25'd541952, -25'd3153175, 25'd1970734}, '{25'd3842932, 25'd1724393, -25'd2512686, 25'd1379514, 25'd2660491, 25'd1872198, 25'd2512686, 25'd492684, -25'd1083904}, '{25'd1280977, 25'd98537, 25'd1921466, 25'd837562, -25'd1428782, 25'd591220, 25'd5173178, 25'd0, 25'd1231709}, '{25'd591220, 25'd2463418, 25'd5567325, -25'd1970734, 25'd197073, 25'd3153175, -25'd1083904, -25'd886830, 25'd1231709}, '{25'd985367, 25'd5518056, 25'd3103907, 25'd3941469, 25'd4631226, 25'd6257082, 25'd4828299, 25'd3793664, -25'd2759028}, '{-25'd1379514, 25'd5468788, 25'd640489, 25'd5370251, 25'd3547322, 25'd5370251, -25'd1625856, 25'd886830, 25'd4926836}, '{25'd591220, -25'd2020003, 25'd3103907, 25'd3202443, -25'd2069271, -25'd2069271, -25'd2857565, 25'd4483421, 25'd197073}, '{25'd2069271, -25'd1872198, -25'd541952, 25'd2217076, -25'd985367, 25'd3744395, -25'd2167808, 25'd3054638, -25'd1724393}}, '{'{25'd640489, -25'd3153175, 25'd1379514, -25'd3005370, 25'd2118539, 25'd2857565, -25'd3793664, 25'd3941469, -25'd2217076}, '{25'd443415, -25'd1478051, -25'd1478051, 25'd3793664, -25'd1527319, 25'd788294, -25'd1379514, -25'd1724393, 25'd443415}, '{25'd3793664, -25'd1527319, -25'd1231709, -25'd1379514, -25'd1478051, -25'd2561955, -25'd1280977, 25'd4335616, -25'd3005370}, '{-25'd4040005, -25'd1724393, -25'd689757, 25'd4040005, 25'd3645859, -25'd3793664, 25'd1724393, 25'd3695127, 25'd0}, '{25'd788294, -25'd739025, 25'd1428782, -25'd2956102, 25'd1773661, 25'd1921466, 25'd788294, 25'd1724393, 25'd2217076}, '{-25'd3596590, 25'd1133172, 25'd2660491, -25'd295610, -25'd344879, 25'd640489, -25'd1083904, -25'd2660491, -25'd837562}, '{25'd2611223, -25'd3941469, 25'd1970734, 25'd5025373, 25'd2709760, 25'd1231709, -25'd1527319, -25'd985367, 25'd3103907}, '{25'd3251712, 25'd98537, 25'd3645859, -25'd936099, 25'd2956102, 25'd4877568, 25'd443415, -25'd2512686, 25'd3744395}, '{25'd2364881, -25'd492684, -25'd1625856, -25'd1182441, -25'd1724393, 25'd4187811, -25'd98537, -25'd1182441, 25'd3842932}}},
    '{'{'{25'd3541958, 25'd715928, -25'd3014432, -25'd904330, 25'd226082, -25'd3843401, 25'd3918762, -25'd1695618, -25'd3052113}, '{25'd3391236, 25'd150722, 25'd1469536, -25'd3730360, 25'd2072422, 25'd3918762, 25'd1431855, 25'd2976752, 25'd1620257}, '{25'd1092732, 25'd2562267, 25'd1205773, 25'd2637628, -25'd3428917, -25'd2863711, 25'd2901391, 25'd527526, 25'd3315875}, '{-25'd904330, 25'd3240515, 25'd3843401, 25'd3014432, -25'd1695618, 25'd2486907, -25'd565206, -25'd753608, -25'd2185463}, '{-25'd904330, -25'd3768040, 25'd339124, 25'd2147783, 25'd2185463, 25'd2449226, 25'd527526, -25'd1884020, 25'd3541958}, '{-25'd3617319, -25'd2260824, -25'd4823092, 25'd3466597, -25'd791288, 25'd1356494, -25'd4069483, -25'd2599948, 25'd1733299}, '{-25'd1770979, -25'd1657938, 25'd2750669, 25'd2373865, 25'd2223144, -25'd3730360, -25'd2712989, -25'd2939071, -25'd3541958}, '{-25'd1620257, 25'd3504277, -25'd4446287, -25'd1507216, 25'd1168092, 25'd2524587, -25'd2939071, -25'd678247, 25'd3654999}, '{25'd3692679, 25'd301443, 25'd3202834, -25'd866649, 25'd2336185, -25'd3278195, -25'd3391236, -25'd2863711, -25'd4107164}}, '{'{-25'd2712989, 25'd226082, -25'd4069483, 25'd1846340, 25'd3994123, 25'd3466597, 25'd1281134, 25'd1356494, 25'd3315875}, '{-25'd678247, -25'd376804, -25'd1808659, 25'd4144844, 25'd1997061, 25'd2336185, -25'd4257885, 25'd2034742, 25'd1921701}, '{25'd1469536, 25'd2788350, 25'd527526, 25'd1846340, -25'd75361, 25'd715928, 25'd1092732, 25'd1921701, -25'd226082}, '{25'd2449226, -25'd2373865, 25'd3843401, 25'd3805721, 25'd791288, -25'd3278195, 25'd791288, -25'd1092732, -25'd1582577}, '{-25'd2486907, 25'd2863711, -25'd1582577, 25'd3617319, 25'd2750669, 25'd1921701, 25'd3843401, -25'd226082, 25'd1997061}, '{25'd3504277, 25'd188402, -25'd4483968, 25'd1808659, 25'd3165154, -25'd2863711, -25'd1092732, 25'd1770979, -25'd828969}, '{-25'd1959381, 25'd1469536, 25'd1168092, -25'd2675309, -25'd753608, 25'd1921701, -25'd1431855, -25'd3353556, -25'd2336185}, '{25'd75361, -25'd2486907, 25'd2185463, 25'd0, -25'd1243453, 25'd565206, 25'd3994123, -25'd2260824, -25'd715928}, '{25'd1846340, 25'd301443, -25'd113041, -25'd791288, 25'd1959381, 25'd1017371, 25'd1959381, 25'd2185463, 25'd1770979}}, '{'{25'd2072422, 25'd1808659, -25'd942010, -25'd1620257, 25'd2599948, 25'd3843401, 25'd1695618, -25'd2147783, -25'd565206}, '{-25'd2901391, -25'd2147783, 25'd1733299, 25'd2223144, 25'd376804, -25'd1318814, -25'd3466597, 25'd4182525, -25'd2939071}, '{25'd4634690, -25'd2373865, -25'd2637628, -25'd1281134, 25'd2147783, 25'd4182525, 25'd3278195, 25'd942010, -25'd3843401}, '{-25'd37680, 25'd4144844, 25'd3768040, 25'd452165, 25'd2486907, 25'd2147783, 25'd3089793, -25'd715928, -25'd904330}, '{25'd4521648, -25'd1997061, -25'd1770979, -25'd3278195, 25'd3504277, -25'd3127473, 25'd452165, 25'd1431855, 25'd1808659}, '{-25'd1997061, -25'd2110103, -25'd414484, -25'd2939071, -25'd3428917, -25'd1733299, 25'd1017371, -25'd1657938, 25'd1997061}, '{-25'd2486907, 25'd2712989, 25'd1921701, 25'd3466597, 25'd2260824, -25'd2976752, 25'd3504277, -25'd1582577, 25'd2034742}, '{25'd2524587, -25'd3617319, -25'd828969, -25'd1243453, 25'd602886, -25'd715928, -25'd1770979, -25'd715928, 25'd1394175}, '{-25'd602886, -25'd4069483, 25'd1884020, -25'd2072422, 25'd489845, 25'd1507216, 25'd678247, -25'd3127473, 25'd263763}}},
    '{'{'{-25'd450384, -25'd2047200, -25'd3357409, 25'd1924368, 25'd3889681, 25'd2333808, 25'd2415697, -25'd450384, 25'd2006256}, '{-25'd4421953, 25'd1514928, 25'd3111745, 25'd859824, 25'd696048, 25'd3029857, 25'd4217233, 25'd40944, 25'd1637760}, '{-25'd777936, -25'd1269264, -25'd1760592, 25'd1064544, 25'd4749505, -25'd3029857, 25'd1392096, 25'd3234577, 25'd696048}, '{-25'd3603073, -25'd5240833, -25'd163776, 25'd3357409, -25'd1473984, 25'd4708561, 25'd3234577, -25'd3521185, -25'd2374753}, '{-25'd4217233, -25'd3029857, -25'd4381009, 25'd1105488, -25'd736992, 25'd3029857, 25'd1392096, -25'd2088144, -25'd573216}, '{-25'd5118001, -25'd2497585, 25'd2497585, -25'd818880, -25'd1637760, 25'd4749505, -25'd1064544, 25'd2702305, -25'd2047200}, '{25'd3398353, -25'd1596816, -25'd2006256, -25'd3193633, 25'd3562129, -25'd2784193, 25'd3725905, 25'd777936, -25'd122832}, '{25'd2947969, -25'd5240833, 25'd1678704, 25'd941712, 25'd1555872, 25'd2170032, 25'd2292864, 25'd1965312, -25'd3562129}, '{-25'd1883424, -25'd368496, -25'd818880, 25'd4217233, 25'd3111745, -25'd3521185, 25'd696048, 25'd2579473, 25'd736992}}, '{'{-25'd2743249, -25'd2579473, -25'd3193633, 25'd1842480, -25'd1883424, 25'd3603073, -25'd1392096, 25'd2866081, -25'd1801536}, '{25'd122832, -25'd4462897, 25'd2210976, 25'd1310208, -25'd2292864, 25'd1555872, 25'd1801536, -25'd2210976, 25'd3234577}, '{-25'd2047200, -25'd2661361, 25'd2210976, 25'd2333808, -25'd818880, 25'd40944, -25'd982656, -25'd1351152, -25'd1801536}, '{-25'd4135345, -25'd777936, -25'd1310208, 25'd2088144, 25'd1555872, -25'd1269264, -25'd2907025, -25'd1801536, -25'd818880}, '{-25'd2988913, -25'd2538529, 25'd3766849, -25'd3684961, -25'd2088144, -25'd982656, 25'd5077057, -25'd40944, -25'd491328}, '{25'd1064544, -25'd4176289, -25'd1801536, -25'd2497585, 25'd1146432, 25'd2579473, -25'd1678704, -25'd1596816, 25'd5118001}, '{-25'd1555872, -25'd2702305, 25'd2497585, 25'd573216, 25'd3480241, 25'd4176289, -25'd2661361, -25'd3029857, -25'd1187376}, '{-25'd573216, -25'd2702305, 25'd1760592, -25'd2415697, -25'd3603073, -25'd900768, -25'd3070801, 25'd2456641, 25'd941712}, '{25'd2907025, -25'd5240833, 25'd163776, 25'd2415697, -25'd3357409, -25'd2743249, -25'd1023600, 25'd2907025, 25'd4217233}}, '{'{-25'd3521185, 25'd2292864, -25'd4135345, -25'd2374753, 25'd2825137, -25'd859824, 25'd1760592, -25'd4544785, -25'd573216}, '{-25'd1064544, -25'd5118001, 25'd163776, -25'd491328, -25'd982656, -25'd4421953, 25'd1760592, 25'd2907025, -25'd2579473}, '{25'd1596816, -25'd4217233, -25'd2988913, 25'd1637760, -25'd1842480, -25'd2907025, 25'd1146432, 25'd3521185, -25'd3275521}, '{25'd3275521, -25'd3971569, -25'd2579473, -25'd2415697, -25'd3889681, 25'd2210976, -25'd327552, -25'd3807793, 25'd3357409}, '{25'd1433040, 25'd3848737, -25'd163776, -25'd3644017, -25'd3111745, -25'd1433040, 25'd368496, -25'd4421953, 25'd655104}, '{25'd409440, -25'd655104, -25'd532272, 25'd1146432, -25'd2538529, -25'd4340065, 25'd2129088, -25'd3766849, -25'd2661361}, '{25'd696048, 25'd3439297, 25'd3193633, 25'd941712, -25'd3930625, -25'd1760592, 25'd3684961, -25'd3398353, 25'd3971569}, '{25'd286608, -25'd2415697, -25'd3357409, 25'd941712, -25'd2579473, -25'd3521185, 25'd3889681, 25'd818880, 25'd2129088}, '{25'd2251920, 25'd2374753, -25'd2292864, 25'd81888, -25'd2210976, -25'd450384, 25'd1678704, 25'd1514928, 25'd368496}}},
    '{'{'{25'd3537087, -25'd1263245, 25'd2737032, 25'd4421359, -25'd589514, -25'd463190, -25'd2484382, -25'd2273842, 25'd3452871}, '{-25'd2315950, -25'd1305353, -25'd2652815, 25'd3663411, -25'd294757, -25'd2821248, 25'd2063301, -25'd1094813, 25'd1052704}, '{25'd4463467, -25'd294757, 25'd463190, 25'd3242330, -25'd3031789, 25'd4295034, -25'd3284438, 25'd4421359, 25'd2821248}, '{25'd5095089, 25'd4295034, 25'd252649, 25'd4716116, -25'd252649, -25'd1094813, 25'd210541, 25'd2989681, -25'd2737032}, '{-25'd1431678, 25'd4716116, -25'd1052704, 25'd2105409, 25'd2484382, -25'd842164, -25'd2947572, -25'd547406, 25'd3873952}, '{-25'd2273842, -25'd3242330, 25'd1389570, -25'd673731, 25'd2105409, -25'd168433, -25'd1810652, -25'd1221137, -25'd2358058}, '{25'd2989681, 25'd1515894, -25'd757947, 25'd2989681, 25'd4126601, -25'd1263245, 25'd42108, -25'd126325, -25'd715839}, '{25'd4126601, 25'd1305353, 25'd1979084, -25'd2568599, -25'd3326546, 25'd4716116, 25'd884272, -25'd757947, 25'd3831844}, '{25'd673731, 25'd1389570, -25'd1389570, 25'd2021192, -25'd3116005, 25'd3747628, -25'd1179029, -25'd505298, 25'd2147517}}, '{'{25'd757947, -25'd3579195, 25'd926380, -25'd2610707, 25'd3116005, -25'd3494979, -25'd1600111, 25'd3116005, -25'd3326546}, '{25'd715839, -25'd4168710, -25'd2021192, -25'd2189625, -25'd4547683, -25'd2105409, 25'd3284438, -25'd1094813, 25'd2737032}, '{-25'd168433, 25'd3452871, -25'd3410762, -25'd3242330, 25'd126325, -25'd3242330, -25'd3368654, 25'd1768543, -25'd2568599}, '{-25'd1179029, -25'd968488, -25'd3831844, -25'd631623, -25'd3916060, 25'd3242330, 25'd3452871, -25'd884272, 25'd2021192}, '{25'd3494979, -25'd673731, 25'd1894868, -25'd5137198, -25'd5221414, -25'd4042385, 25'd2652815, 25'd1136921, -25'd210541}, '{25'd2821248, -25'd4252926, -25'd2484382, -25'd1979084, -25'd4337142, -25'd3789736, 25'd1979084, -25'd3663411, 25'd4589791}, '{25'd1979084, 25'd1558003, -25'd1136921, 25'd294757, -25'd4379250, 25'd463190, 25'd2863356, -25'd2694923, -25'd3073897}, '{25'd884272, -25'd631623, -25'd2442274, -25'd673731, -25'd4210818, -25'd2821248, 25'd336865, 25'd2021192, -25'd3242330}, '{25'd1936976, 25'd547406, -25'd3073897, 25'd3452871, 25'd2021192, 25'd2694923, -25'd3368654, -25'd3116005, -25'd3242330}}, '{'{-25'd3031789, 25'd3958169, 25'd378974, 25'd4126601, -25'd1810652, 25'd3242330, 25'd1094813, 25'd252649, 25'd2526491}, '{25'd3284438, -25'd2442274, 25'd2863356, -25'd1810652, 25'd3789736, -25'd505298, 25'd5221414, 25'd5052981, -25'd1684327}, '{-25'd3200221, 25'd4716116, 25'd2652815, 25'd5263522, 25'd1515894, -25'd3494979, 25'd2905464, -25'd3116005, 25'd2652815}, '{25'd4000277, 25'd84216, 25'd4084493, 25'd800055, 25'd3242330, 25'd3073897, 25'd1515894, -25'd673731, 25'd2652815}, '{-25'd1052704, -25'd2273842, 25'd2652815, 25'd1642219, 25'd3410762, 25'd1894868, 25'd1558003, 25'd1894868, 25'd4968765}, '{25'd757947, 25'd1347462, 25'd3073897, -25'd2863356, -25'd3326546, -25'd1810652, -25'd3452871, -25'd1136921, 25'd463190}, '{-25'd378974, 25'd2189625, 25'd3789736, -25'd252649, 25'd4631899, -25'd1768543, -25'd1263245, -25'd1768543, 25'd673731}, '{25'd715839, 25'd5347738, -25'd715839, 25'd2442274, -25'd3031789, -25'd968488, 25'd3073897, 25'd1179029, 25'd4000277}, '{25'd3116005, 25'd3284438, 25'd2947572, -25'd2652815, 25'd2021192, 25'd4589791, -25'd84216, 25'd2021192, 25'd1726435}}},
    '{'{'{-25'd543838, 25'd4241938, -25'd4350705, 25'd2429144, 25'd2791703, 25'd1341468, -25'd1196444, -25'd2429144, 25'd145024}, '{-25'd3661844, -25'd2284120, 25'd833885, -25'd2139097, -25'd3879379, 25'd4350705, 25'd1921562, -25'd1994073, 25'd398815}, '{-25'd3190517, 25'd543838, -25'd290047, 25'd870141, -25'd1305212, 25'd108768, 25'd36256, 25'd217535, -25'd507582}, '{25'd4314450, 25'd2936726, -25'd36256, 25'd725118, 25'd761373, -25'd3480564, -25'd1413979, -25'd1812794, -25'd2066585}, '{-25'd3299285, 25'd3335541, 25'd4169426, -25'd3118006, 25'd4350705, 25'd1196444, 25'd507582, -25'd3625588, -25'd398815}, '{25'd2465400, 25'd3371797, -25'd870141, -25'd2284120, 25'd1160188, -25'd2574167, 25'd2211609, -25'd2392888, 25'd616350}, '{25'd1522747, -25'd1667770, -25'd435071, -25'd1667770, -25'd4060658, 25'd0, 25'd1341468, -25'd4060658, 25'd1015165}, '{25'd1957817, 25'd2139097, -25'd761373, 25'd833885, -25'd2175353, 25'd253791, -25'd3081750, 25'd2320376, 25'd145024}, '{-25'd108768, 25'd2610423, 25'd253791, -25'd833885, -25'd253791, 25'd1160188, -25'd3734355, 25'd1087676, 25'd4169426}}, '{'{25'd0, 25'd1015165, -25'd2211609, 25'd507582, -25'd362559, 25'd3516820, -25'd1994073, -25'd1704026, 25'd3154261}, '{25'd652606, 25'd1957817, -25'd3045494, 25'd2972982, 25'd2501656, -25'd3154261, 25'd4133170, -25'd362559, 25'd797629}, '{-25'd435071, -25'd1015165, -25'd1885306, -25'd3480564, -25'd4096914, 25'd2972982, 25'd1051420, -25'd2900470, 25'd4241938}, '{-25'd1123932, -25'd1631515, -25'd362559, -25'd3770611, 25'd797629, 25'd3045494, 25'd1595259, -25'd4060658, -25'd2574167}, '{-25'd1486491, 25'd688862, -25'd797629, 25'd3879379, -25'd1196444, -25'd4096914, -25'd471326, 25'd2827959, -25'd3444308}, '{25'd3843123, -25'd2356632, 25'd906397, 25'd3516820, 25'd1160188, 25'd1341468, 25'd3553076, -25'd2646679, 25'd942653}, '{25'd2719191, 25'd3226773, 25'd1704026, 25'd2211609, -25'd1522747, 25'd3045494, 25'd2537911, -25'd2537911, 25'd978909}, '{25'd2501656, 25'd2972982, 25'd2755447, -25'd2211609, 25'd3843123, -25'd978909, -25'd4241938, -25'd2900470, 25'd906397}, '{-25'd3190517, -25'd435071, -25'd72512, -25'd652606, -25'd2356632, -25'd543838, 25'd3734355, 25'd652606, -25'd725118}}, '{'{-25'd2247864, -25'd2719191, 25'd3951891, -25'd580094, 25'd2211609, -25'd3226773, -25'd3154261, -25'd181279, -25'd1123932}, '{-25'd1776538, -25'd1885306, -25'd2574167, 25'd2356632, 25'd3625588, 25'd2719191, 25'd4350705, -25'd2066585, -25'd1631515}, '{-25'd3951891, -25'd4205682, 25'd870141, 25'd1051420, 25'd2320376, 25'd2501656, 25'd507582, -25'd3154261, -25'd2139097}, '{25'd2900470, -25'd3770611, 25'd145024, 25'd4531985, 25'd2465400, 25'd3698100, 25'd725118, -25'd2574167, 25'd362559}, '{-25'd4133170, 25'd2864214, -25'd1413979, 25'd2682935, -25'd1667770, 25'd2465400, 25'd4604497, -25'd1776538, 25'd978909}, '{-25'd2175353, 25'd2936726, -25'd1232700, -25'd1305212, -25'd3480564, 25'd3371797, 25'd4604497, 25'd2574167, -25'd942653}, '{-25'd1196444, -25'd2392888, 25'd145024, 25'd3408053, 25'd2610423, -25'd3661844, 25'd4096914, 25'd1812794, 25'd3444308}, '{25'd181279, 25'd3335541, 25'd797629, -25'd3226773, 25'd4350705, 25'd1160188, -25'd2646679, 25'd543838, 25'd1885306}, '{-25'd2610423, 25'd1849050, 25'd3951891, 25'd543838, 25'd1305212, 25'd1087676, 25'd3553076, 25'd2465400, -25'd4060658}}},
    '{'{'{25'd2036020, -25'd2639285, -25'd980306, 25'd2865509, -25'd377041, 25'd1319642, -25'd1357347, 25'd4072040, 25'd2224540}, '{25'd4147448, -25'd2149132, 25'd1885204, -25'd4147448, 25'd829490, -25'd3054030, 25'd3544183, -25'd377041, 25'd3845815}, '{25'd2036020, 25'd3770407, -25'd2790101, 25'd490153, 25'd1018010, -25'd2036020, -25'd4185152, -25'd188520, 25'd2752397}, '{-25'd1357347, -25'd3317958, 25'd2827805, -25'd4260560, -25'd2111428, 25'd2111428, 25'd3280254, -25'd1131122, -25'd1470459}, '{-25'd716377, 25'd980306, -25'd4335968, -25'd1206530, 25'd1508163, -25'd2375356, -25'd4411376, 25'd1395051, 25'd1470459}, '{25'd3506479, 25'd490153, 25'd1658979, 25'd565561, -25'd3355662, -25'd377041, 25'd2337652, -25'd1508163, -25'd1206530}, '{25'd1432755, -25'd904898, -25'd1357347, -25'd3921223, -25'd339337, -25'd3431070, 25'd339337, 25'd2903213, -25'd2337652}, '{-25'd829490, -25'd1018010, 25'd678673, -25'd1206530, 25'd3732703, -25'd3054030, 25'd2488469, 25'd640969, -25'd603265}, '{25'd3468775, -25'd3845815, 25'd2601581, 25'd2752397, -25'd3996632, -25'd3242550, -25'd1055714, 25'd1809795, 25'd3694999}}, '{'{-25'd1922908, -25'd2526173, 25'd113112, 25'd4298264, 25'd1319642, 25'd1545867, 25'd1847499, 25'd565561, -25'd867194}, '{25'd3619591, 25'd2149132, -25'd2601581, 25'd2563877, -25'd3393366, -25'd2940918, -25'd1545867, -25'd3091734, -25'd3845815}, '{25'd3431070, 25'd1470459, -25'd2903213, -25'd3732703, -25'd4222856, -25'd2186836, 25'd2978622, -25'd3770407, 25'd4109744}, '{-25'd603265, -25'd3694999, -25'd2827805, 25'd1395051, -25'd2526173, -25'd3317958, 25'd3506479, -25'd1696683, -25'd1357347}, '{25'd2036020, 25'd4449080, 25'd1244234, 25'd339337, -25'd527857, 25'd1244234, 25'd2149132, 25'd377041, -25'd2488469}, '{-25'd829490, 25'd3619591, 25'd1093418, 25'd1055714, 25'd3317958, -25'd4373672, 25'd1696683, -25'd339337, 25'd942602}, '{-25'd3129438, -25'd3431070, -25'd3581887, 25'd4222856, 25'd2940918, -25'd2337652, -25'd2714693, -25'd2186836, -25'd1696683}, '{-25'd1093418, -25'd1131122, -25'd3393366, -25'd1432755, -25'd1281938, 25'd1847499, 25'd3619591, 25'd1470459, 25'd4675305}, '{25'd1319642, 25'd4373672, -25'd603265, 25'd4298264, -25'd339337, 25'd414745, 25'd1395051, 25'd4713009, -25'd1206530}}, '{'{25'd3732703, -25'd75408, -25'd1960612, -25'd3958927, -25'd2865509, 25'd3694999, -25'd3054030, 25'd2299948, -25'd3204846}, '{25'd640969, 25'd4034336, -25'd1093418, -25'd2903213, 25'd1432755, 25'd1658979, -25'd2865509, 25'd867194, -25'd490153}, '{-25'd2827805, 25'd1508163, 25'd2714693, 25'd1545867, -25'd603265, -25'd904898, -25'd2676989, 25'd3468775, 25'd3129438}, '{-25'd980306, 25'd678673, 25'd2865509, -25'd678673, -25'd3694999, -25'd2827805, -25'd3958927, -25'd1018010, 25'd4373672}, '{25'd1960612, 25'd150816, -25'd1168826, -25'd4072040, 25'd3544183, -25'd2827805, -25'd3468775, -25'd1847499, 25'd2111428}, '{-25'd2111428, 25'd3544183, 25'd2111428, -25'd942602, -25'd339337, 25'd1960612, -25'd1998316, -25'd1319642, 25'd226224}, '{-25'd3770407, 25'd4788417, 25'd904898, 25'd2752397, 25'd1847499, -25'd1470459, 25'd3694999, -25'd1658979, -25'd1093418}, '{25'd301633, -25'd942602, 25'd942602, -25'd3167142, -25'd1319642, 25'd1206530, 25'd1470459, -25'd2149132, 25'd452449}, '{-25'd3581887, 25'd3317958, -25'd188520, -25'd3431070, 25'd2714693, 25'd3845815, 25'd1696683, 25'd1847499, 25'd3317958}}},
    '{'{'{-25'd1771286, -25'd3072639, 25'd4518587, 25'd4446289, -25'd1988178, 25'd3036490, -25'd2096624, -25'd2530409, 25'd1662840}, '{25'd3253382, -25'd3289531, 25'd2205070, 25'd2964193, 25'd1409799, -25'd614528, 25'd1482096, 25'd3904059, 25'd2783449}, '{25'd1337502, 25'd4554735, -25'd2891895, 25'd3361828, 25'd1156758, -25'd903717, -25'd1301353, 25'd1048312, 25'd3181085}, '{25'd1735137, 25'd4193248, -25'd2385814, -25'd903717, -25'd2928044, -25'd1952029, 25'd831420, 25'd108446, 25'd2241219}, '{-25'd3651018, 25'd4590884, -25'd3470275, -25'd36149, -25'd1771286, 25'd108446, -25'd36149, -25'd3651018, -25'd3687167}, '{25'd759123, 25'd3181085, -25'd1084461, -25'd2458111, -25'd2132773, -25'd2385814, -25'd469933, 25'd469933, -25'd1518245}, '{-25'd72297, 25'd722974, -25'd144595, -25'd108446, 25'd4120951, 25'd180743, 25'd542230, 25'd3795613, 25'd2060476}, '{-25'd4012505, -25'd2205070, 25'd3614869, 25'd397636, -25'd1192907, 25'd1445948, 25'd4084802, 25'd2421962, 25'd2747301}, '{25'd2747301, -25'd1590543, 25'd2891895, 25'd1265204, -25'd72297, -25'd3397977, 25'd1662840, 25'd3434126, -25'd361487}}, '{'{-25'd2891895, 25'd1735137, 25'd831420, -25'd3253382, -25'd3904059, -25'd3181085, -25'd1518245, 25'd1337502, 25'd2096624}, '{-25'd1409799, 25'd2060476, -25'd2711152, -25'd4084802, 25'd2494260, -25'd361487, -25'd1120609, -25'd3542572, -25'd2349665}, '{-25'd3831762, -25'd3542572, 25'd2638855, -25'd1084461, 25'd361487, -25'd1518245, 25'd3651018, 25'd1012163, 25'd2132773}, '{25'd3867910, 25'd2385814, 25'd2638855, -25'd361487, -25'd3397977, 25'd1735137, 25'd1012163, -25'd289190, 25'd2855747}, '{-25'd2530409, -25'd3651018, 25'd3470275, -25'd2421962, 25'd1735137, -25'd433784, 25'd3470275, 25'd1156758, -25'd3723315}, '{-25'd2747301, -25'd578379, -25'd1554394, -25'd578379, 25'd3434126, 25'd325338, 25'd2349665, -25'd3723315, -25'd686825}, '{25'd2638855, -25'd2385814, 25'd3759464, -25'd3976356, 25'd2855747, -25'd650676, 25'd1735137, 25'd1084461, -25'd1771286}, '{25'd506082, -25'd3217234, -25'd3976356, -25'd1156758, -25'd3795613, -25'd614528, -25'd1879732, -25'd3578721, -25'd144595}, '{25'd180743, 25'd831420, 25'd2675003, 25'd72297, -25'd361487, -25'd3506423, 25'd4590884, 25'd216892, -25'd1554394}}, '{'{25'd3542572, 25'd1554394, -25'd3867910, -25'd2060476, -25'd939866, -25'd2819598, 25'd3687167, -25'd2602706, 25'd1337502}, '{-25'd2385814, -25'd1048312, -25'd976015, 25'd1301353, 25'd2168922, 25'd1229056, 25'd3434126, 25'd3072639, 25'd1807435}, '{-25'd795271, -25'd3108788, -25'd2096624, -25'd144595, -25'd3976356, 25'd2783449, -25'd289190, -25'd1626691, -25'd1735137}, '{-25'd2494260, 25'd4337843, 25'd4301695, -25'd3361828, 25'd2928044, 25'd1879732, 25'd3470275, 25'd3723315, -25'd397636}, '{25'd3687167, -25'd2819598, -25'd72297, -25'd3072639, 25'd4590884, 25'd2928044, 25'd3976356, 25'd3325680, 25'd3470275}, '{25'd1590543, 25'd3867910, 25'd1662840, 25'd3651018, -25'd2928044, 25'd939866, 25'd3506423, 25'd2566557, -25'd1156758}, '{25'd4301695, 25'd3651018, -25'd253041, 25'd2566557, 25'd867569, 25'd2964193, -25'd1807435, -25'd3723315, 25'd3434126}, '{25'd180743, -25'd3181085, -25'd2421962, 25'd216892, -25'd2964193, -25'd2964193, 25'd4482438, 25'd867569, 25'd2819598}, '{-25'd2928044, -25'd3397977, -25'd3614869, 25'd216892, -25'd3904059, -25'd1843583, -25'd650676, 25'd4120951, 25'd1698989}}},
    '{'{'{-25'd4188334, -25'd1754089, -25'd2935414, 25'd751752, 25'd3937750, 25'd2291055, 25'd680157, 25'd894943, 25'd2935414}, '{25'd393775, -25'd1038134, 25'd3722964, 25'd1324516, -25'd1360314, 25'd3508178, 25'd608561, -25'd1503505, -25'd536966}, '{25'd3114403, -25'd3937750, 25'd1038134, -25'd3866155, 25'd787550, -25'd1145527, -25'd2112066, -25'd1861482, 25'd3722964}, '{25'd608561, -25'd1897280, 25'd2219459, -25'd4116739, -25'd107393, 25'd2326852, -25'd3436582, 25'd178989, 25'd680157}, '{25'd2147864, -25'd1825684, -25'd751752, 25'd2828021, -25'd2040471, -25'd178989, 25'd71595, -25'd3472380, -25'd3937750}, '{25'd608561, -25'd3937750, -25'd3114403, -25'd2076268, 25'd2971212, 25'd3472380, 25'd3436582, -25'd787550, 25'd1073932}, '{-25'd2434246, 25'd1575100, -25'd2649032, 25'd1002336, 25'd4116739, 25'd393775, -25'd3937750, -25'd3293391, -25'd2147864}, '{-25'd35798, -25'd1360314, -25'd1109730, 25'd322180, 25'd4080941, 25'd465370, -25'd3221796, 25'd3400784, -25'd966539}, '{25'd178989, 25'd536966, -25'd2183662, -25'd3508178, 25'd4116739, 25'd1503505, 25'd1467707, 25'd4438919, -25'd3185998}}, '{'{-25'd71595, -25'd1360314, 25'd4438919, -25'd751752, 25'd2649032, 25'd3794559, 25'd1789887, 25'd1109730, 25'd859146}, '{25'd3579773, 25'd4259930, -25'd3293391, 25'd2470043, 25'd143191, 25'd4546312, 25'd2040471, -25'd2470043, -25'd4045143}, '{25'd4259930, -25'd1610898, 25'd966539, 25'd751752, 25'd3150200, -25'd3901953, 25'd1288718, 25'd572764, 25'd2040471}, '{25'd2541639, 25'd644359, 25'd751752, -25'd3758762, 25'd2649032, -25'd1503505, -25'd1754089, 25'd3042807, 25'd1145527}, '{-25'd715955, 25'd1109730, -25'd1288718, -25'd2255257, 25'd4259930, -25'd250584, 25'd3293391, -25'd3472380, -25'd1968875}, '{25'd1539302, 25'd1861482, 25'd4295728, -25'd4259930, -25'd2649032, -25'd2147864, -25'd1646696, 25'd715955, -25'd2112066}, '{-25'd2935414, -25'd1825684, 25'd2326852, 25'd3221796, -25'd2291055, -25'd3758762, -25'd3364987, -25'd4045143, 25'd2255257}, '{25'd1646696, -25'd3830357, -25'd2434246, -25'd322180, 25'd3329189, 25'd1575100, -25'd2362650, -25'd572764, 25'd3078605}, '{25'd644359, -25'd3687166, 25'd894943, 25'd787550, 25'd1861482, -25'd3651368, 25'd1933077, 25'd2971212, 25'd4295728}}, '{'{-25'd214786, -25'd2649032, -25'd71595, -25'd572764, -25'd3293391, 25'd4080941, -25'd1968875, 25'd465370, 25'd2326852}, '{-25'd3150200, 25'd1861482, 25'd107393, -25'd787550, 25'd4510514, 25'd966539, 25'd4438919, -25'd1181325, -25'd2756425}, '{25'd4438919, 25'd3830357, -25'd1968875, 25'd2147864, -25'd2577437, -25'd3830357, 25'd1431909, 25'd3150200, 25'd4259930}, '{-25'd1396111, -25'd1897280, -25'd2362650, -25'd2899616, -25'd1217123, 25'd2684830, -25'd2112066, -25'd572764, -25'd4224132}, '{25'd3722964, 25'd3758762, 25'd2577437, -25'd644359, -25'd3508178, 25'd4080941, -25'd4367323, -25'd3007009, -25'd3185998}, '{25'd286382, -25'd2684830, -25'd322180, -25'd3579773, 25'd3293391, -25'd4045143, 25'd2505841, -25'd2326852, -25'd3400784}, '{25'd2398448, 25'd1109730, 25'd3078605, 25'd250584, 25'd2613234, 25'd4009346, -25'd3901953, -25'd1252921, -25'd1217123}, '{25'd3794559, 25'd966539, 25'd1754089, 25'd3937750, -25'd1503505, 25'd3078605, 25'd1610898, 25'd2720627, -25'd1431909}, '{25'd2828021, -25'd3579773, -25'd2040471, -25'd4080941, -25'd71595, -25'd1539302, 25'd4116739, -25'd536966, 25'd3150200}}},
    '{'{'{25'd468385, 25'd2877221, 25'd5352969, -25'd1672803, -25'd2743396, -25'd4817672, 25'd1338242, 25'd334561, 25'd802945}, '{-25'd4416199, -25'd869857, 25'd5620617, 25'd2609572, 25'd1605891, -25'd535297, 25'd267648, 25'd200736, 25'd267648}, '{25'd2743396, 25'd4215463, 25'd602209, -25'd736033, -25'd2208100, -25'd4550023, -25'd4215463, -25'd535297, -25'd66912}, '{25'd5352969, 25'd3011045, 25'd4483111, 25'd3747078, -25'd2810309, -25'd1605891, -25'd3613254, -25'd6089002, 25'd869857}, '{25'd133824, 25'd3546342, 25'd5018408, -25'd1204418, -25'd7293420, -25'd4550023, -25'd5687529, -25'd2141187, -25'd2676484}, '{25'd1472066, 25'd2542660, 25'd3880902, -25'd2877221, -25'd2475748, -25'd2542660, -25'd6624299, 25'd3278693, 25'd6423562}, '{25'd4483111, 25'd602209, 25'd4951496, 25'd1538978, -25'd2208100, 25'd2676484, -25'd3813990, 25'd3813990, 25'd4215463}, '{-25'd5018408, 25'd2676484, -25'd3613254, -25'd3880902, 25'd1204418, -25'd2676484, -25'd5286057, -25'd4616935, -25'd2475748}, '{-25'd3077957, -25'd6490475, -25'd1538978, -25'd401473, 25'd2542660, 25'd3813990, 25'd7025771, -25'd1940451, -25'd1472066}}, '{'{25'd802945, 25'd3479430, -25'd936770, 25'd602209, 25'd2877221, -25'd1003682, 25'd200736, -25'd6691211, -25'd936770}, '{25'd2877221, -25'd1873539, -25'd1338242, 25'd5486793, 25'd535297, 25'd3613254, 25'd1137506, 25'd2609572, 25'd3747078}, '{25'd4884584, 25'd1271330, 25'd5219144, 25'd2208100, -25'd2877221, -25'd267648, 25'd2141187, -25'd66912, -25'd4550023}, '{25'd2141187, 25'd535297, 25'd5687529, -25'd2877221, -25'd736033, -25'd4750760, -25'd5888266, -25'd66912, -25'd1405154}, '{25'd2074275, 25'd4616935, 25'd5888266, 25'd1070594, 25'd1137506, 25'd0, -25'd5687529, -25'd6155914, -25'd2944133}, '{25'd3680166, 25'd8497838, 25'd2743396, 25'd1137506, 25'd736033, -25'd2810309, 25'd1472066, -25'd4951496, 25'd3412518}, '{25'd6958859, 25'd468385, -25'd602209, -25'd3144869, 25'd2275012, -25'd2810309, -25'd736033, -25'd2676484, 25'd1137506}, '{-25'd4483111, 25'd3077957, -25'd2141187, -25'd2542660, -25'd3278693, 25'd3880902, -25'd1605891, -25'd7962541, -25'd3813990}, '{25'd401473, 25'd2542660, -25'd2542660, 25'd1338242, 25'd1739715, 25'd2475748, 25'd4215463, -25'd2475748, -25'd6490475}}, '{'{-25'd6423562, -25'd3077957, -25'd4416199, -25'd3345605, -25'd1472066, 25'd669121, -25'd1605891, -25'd535297, 25'd1405154}, '{-25'd4750760, -25'd4483111, 25'd401473, 25'd4081639, -25'd3345605, -25'd3345605, -25'd3747078, -25'd1538978, 25'd2877221}, '{-25'd334561, 25'd4951496, 25'd936770, -25'd669121, 25'd3412518, -25'd1070594, -25'd2676484, -25'd200736, 25'd936770}, '{-25'd535297, 25'd5286057, 25'd4951496, -25'd669121, 25'd1873539, 25'd2074275, -25'd4148551, -25'd4215463, 25'd7092684}, '{25'd4817672, 25'd3412518, 25'd5620617, 25'd5553705, -25'd3345605, -25'd869857, -25'd3947814, -25'd802945, 25'd4550023}, '{25'd1338242, 25'd3680166, 25'd1538978, 25'd3747078, 25'd736033, -25'd8364014, -25'd468385, 25'd133824, 25'd3479430}, '{-25'd869857, 25'd4951496, -25'd936770, 25'd3412518, -25'd6022090, 25'd0, -25'd5018408, -25'd4750760, 25'd3479430}, '{-25'd3011045, 25'd200736, 25'd1940451, -25'd2141187, -25'd2877221, -25'd3613254, -25'd736033, -25'd2275012, -25'd3813990}, '{-25'd2944133, -25'd5219144, -25'd3947814, 25'd1271330, 25'd535297, 25'd4750760, 25'd2141187, 25'd1940451, 25'd4750760}}},
    '{'{'{-25'd435306, -25'd72551, 25'd2103977, -25'd181377, 25'd3736374, 25'd3301068, -25'd2829487, 25'd1487294, -25'd2140253}, '{-25'd1704947, -25'd2140253, 25'd4207955, 25'd906887, 25'd4280506, -25'd834336, 25'd1668672, 25'd36275, -25'd2503008}, '{-25'd616683, 25'd1632396, 25'd1414743, 25'd4389332, 25'd652959, 25'd1886325, -25'd2974589, 25'd362755, -25'd2829487}, '{25'd4062853, -25'd689234, -25'd2430457, -25'd1051989, 25'd1777498, -25'd2103977, -25'd108826, -25'd3409895, 25'd3228517}, '{-25'd1160815, -25'd2648110, 25'd2575559, -25'd2466732, -25'd616683, 25'd1850049, -25'd1269642, -25'd3264793, 25'd870611}, '{-25'd1051989, 25'd2575559, -25'd72551, 25'd4171679, -25'd2103977, -25'd3518721, 25'd1088264, -25'd217653, 25'd834336}, '{-25'd399030, -25'd725509, -25'd3228517, 25'd4171679, 25'd3917751, -25'd1704947, -25'd471581, -25'd1197091, 25'd1414743}, '{25'd1305917, 25'd3264793, 25'd4171679, 25'd2865762, -25'd3301068, 25'd616683, -25'd1160815, 25'd1378468, 25'd1451019}, '{25'd2938313, 25'd2829487, -25'd2103977, 25'd544132, 25'd3083415, -25'd1487294, 25'd4244230, -25'd1704947, 25'd399030}}, '{'{-25'd4099128, -25'd725509, -25'd3772649, -25'd3772649, 25'd2974589, 25'd4570710, -25'd2394181, 25'd906887, 25'd4099128}, '{25'd3700098, 25'd3990302, 25'd725509, -25'd761785, -25'd3482445, -25'd145102, 25'd72551, -25'd2466732, 25'd798060}, '{25'd3373619, 25'd2611834, 25'd2902038, 25'd2974589, -25'd2575559, -25'd2793211, 25'd3736374, -25'd2249079, 25'd4135404}, '{25'd4280506, -25'd1922600, -25'd1922600, 25'd3917751, 25'd2430457, 25'd3881476, 25'd72551, 25'd3228517, 25'd1124540}, '{25'd36275, 25'd2829487, 25'd652959, 25'd1632396, -25'd326479, 25'd3155966, 25'd2720661, -25'd2938313, 25'd181377}, '{25'd1958876, 25'd362755, 25'd4353057, -25'd1233366, -25'd3845200, 25'd2466732, -25'd1632396, -25'd1632396, -25'd2176528}, '{-25'd3373619, -25'd3808925, -25'd1958876, 25'd1342193, -25'd1886325, -25'd36275, 25'd1850049, 25'd4606985, -25'd2285355}, '{-25'd689234, 25'd3482445, -25'd3881476, 25'd1850049, 25'd1305917, -25'd2648110, -25'd2249079, -25'd870611, -25'd1704947}, '{25'd3228517, 25'd1850049, -25'd3954027, -25'd2212804, -25'd3337344, 25'd181377, -25'd834336, 25'd1051989, 25'd2539283}}, '{'{25'd4207955, -25'd1886325, -25'd1378468, -25'd2249079, 25'd3409895, -25'd1777498, 25'd4171679, 25'd4316781, 25'd1269642}, '{25'd3772649, 25'd2902038, -25'd3373619, -25'd108826, -25'd3845200, -25'd2974589, 25'd2756936, -25'd689234, -25'd1269642}, '{25'd3010864, -25'd1559845, -25'd290204, 25'd943162, 25'd2430457, 25'd761785, -25'd3808925, 25'd1233366, 25'd3119691}, '{-25'd2648110, 25'd290204, -25'd943162, -25'd2357906, -25'd2974589, -25'd1777498, 25'd4135404, -25'd3409895, 25'd2902038}, '{25'd652959, -25'd1995151, -25'd4171679, 25'd2140253, -25'd2212804, 25'd616683, 25'd3808925, -25'd1632396, -25'd1414743}, '{-25'd3482445, -25'd1414743, -25'd1777498, 25'd3337344, -25'd2575559, 25'd217653, 25'd580408, 25'd2103977, -25'd217653}, '{25'd3083415, 25'd2394181, -25'd3228517, -25'd1596121, 25'd689234, -25'd2756936, 25'd3119691, -25'd4135404, -25'd326479}, '{-25'd471581, -25'd3700098, 25'd761785, 25'd507857, -25'd2938313, -25'd3047140, -25'd3736374, 25'd3518721, -25'd3990302}, '{25'd2103977, 25'd1160815, -25'd3409895, 25'd3954027, 25'd3808925, 25'd399030, 25'd834336, 25'd3119691, 25'd3990302}}},
    '{'{'{25'd1171366, 25'd0, -25'd5135989, -25'd90105, -25'd270315, -25'd5766725, -25'd4730516, 25'd2477890, -25'd4865674}, '{-25'd3333888, 25'd3694308, -25'd1937259, 25'd4279991, -25'd1531786, -25'd1757049, -25'd1982312, -25'd4234938, -25'd4460201}, '{25'd2162522, 25'd1126313, 25'd180210, 25'd2838310, 25'd4640411, -25'd3649255, 25'd0, -25'd1441681, -25'd2613047}, '{-25'd3018520, -25'd3649255, 25'd2207574, -25'd1081261, 25'd2072417, -25'd180210, 25'd2207574, 25'd3469045, -25'd2207574}, '{25'd180210, -25'd2252627, 25'd2117469, 25'd2072417, 25'd4279991, -25'd2297679, -25'd2928415, 25'd3784413, 25'd765893}, '{25'd3063572, 25'd1261471, -25'd315368, 25'd2387784, 25'd3378940, -25'd3018520, -25'd1396629, 25'd2117469, 25'd2432837}, '{25'd1306524, 25'd450525, 25'd3604203, 25'd3514098, 25'd405473, 25'd360420, 25'd1216418, 25'd3063572, 25'd630736}, '{-25'd1576839, 25'd1621891, -25'd360420, -25'd270315, -25'd495578, 25'd2883362, -25'd2117469, -25'd1306524, 25'd1757049}, '{-25'd2207574, 25'd2973467, -25'd810946, -25'd3288835, 25'd4640411, -25'd3378940, 25'd3694308, -25'd3694308, -25'd1036208}}, '{'{-25'd4595359, -25'd901051, -25'd1261471, 25'd360420, -25'd4550306, -25'd360420, -25'd1486734, -25'd4370096, 25'd3469045}, '{25'd2252627, 25'd2883362, -25'd45053, 25'd3378940, 25'd991156, -25'd810946, -25'd495578, -25'd1036208, -25'd3784413}, '{25'd2117469, 25'd3288835, 25'd675788, -25'd1621891, 25'd3604203, 25'd225263, -25'd4325043, -25'd3559150, 25'd3333888}, '{-25'd3739361, 25'd540630, 25'd2387784, 25'd450525, 25'd901051, -25'd3919571, 25'd180210, 25'd3333888, -25'd3423993}, '{-25'd2162522, 25'd765893, 25'd1937259, 25'd3829466, 25'd4279991, -25'd540630, 25'd1531786, -25'd2162522, -25'd4189886}, '{-25'd1757049, 25'd3018520, -25'd225263, -25'd1126313, -25'd270315, -25'd1351576, 25'd135158, 25'd2883362, -25'd1396629}, '{25'd90105, -25'd4144833, 25'd1531786, -25'd765893, 25'd2658100, 25'd225263, -25'd3559150, 25'd315368, 25'd991156}, '{25'd675788, -25'd4595359, 25'd1441681, 25'd901051, -25'd1847154, -25'd1576839, -25'd1216418, 25'd2522942, -25'd4325043}, '{25'd1351576, -25'd495578, 25'd630736, 25'd3739361, 25'd4415149, -25'd1306524, 25'd810946, 25'd3423993, -25'd4685464}}, '{'{25'd180210, -25'd2567995, -25'd810946, -25'd1757049, -25'd3694308, -25'd5045884, -25'd2297679, 25'd4325043, 25'd2432837}, '{-25'd135158, 25'd3559150, 25'd3964623, 25'd3108625, 25'd991156, 25'd1351576, -25'd1847154, 25'd4730516, -25'd360420}, '{-25'd1081261, 25'd1171366, 25'd946103, -25'd1261471, 25'd2162522, -25'd810946, -25'd1847154, -25'd675788, 25'd4009676}, '{25'd1396629, -25'd1757049, 25'd2793257, 25'd3829466, -25'd1261471, -25'd675788, 25'd1802101, -25'd3018520, -25'd315368}, '{-25'd4189886, -25'd3784413, 25'd2432837, -25'd2432837, 25'd3333888, -25'd2883362, 25'd1621891, -25'd2522942, 25'd0}, '{25'd2162522, -25'd1531786, 25'd450525, -25'd1171366, 25'd2522942, 25'd3829466, -25'd991156, 25'd3874518, 25'd2117469}, '{-25'd3423993, -25'd3784413, -25'd946103, 25'd2477890, 25'd4820621, -25'd495578, -25'd3198730, -25'd2477890, -25'd2477890}, '{-25'd3243783, -25'd2162522, -25'd855998, 25'd1802101, 25'd3469045, 25'd1982312, 25'd4550306, -25'd2477890, -25'd225263}, '{-25'd4189886, 25'd180210, 25'd1982312, -25'd3198730, 25'd855998, -25'd1306524, 25'd630736, -25'd3018520, -25'd1036208}}},
    '{'{'{25'd3858640, -25'd2778221, 25'd4514609, -25'd655969, 25'd4051572, 25'd1582042, -25'd3009739, -25'd3434189, 25'd2430943}, '{25'd2623875, 25'd4244504, 25'd3897226, 25'd308691, 25'd115759, 25'd4090158, 25'd3704294, 25'd771728, -25'd1041833}, '{-25'd2508116, -25'd578796, 25'd192932, 25'd231518, 25'd1582042, 25'd2662461, 25'd926074, -25'd347278, 25'd1311938}, '{25'd1273351, 25'd231518, 25'd347278, -25'd2045079, -25'd1620629, 25'd1659215, -25'd501623, -25'd655969, 25'd3588535}, '{25'd4283090, 25'd270105, -25'd655969, 25'd3511362, -25'd1350524, 25'd192932, 25'd2932566, -25'd4090158, 25'd1157592}, '{25'd192932, 25'd1543456, -25'd1119006, -25'd1196178, 25'd1543456, -25'd3048325, 25'd4167331, 25'd3627121, 25'd1774974}, '{-25'd4051572, -25'd2045079, -25'd2238011, -25'd1234765, -25'd2855393, 25'd2469529, 25'd2778221, 25'd4514609, -25'd3897226}, '{25'd1504870, -25'd3279844, 25'd2430943, 25'd2122252, 25'd115759, -25'd810314, -25'd1389110, -25'd2006493, -25'd2238011}, '{25'd1196178, -25'd655969, 25'd2508116, 25'd578796, 25'd2739634, -25'd3125498, 25'd38586, 25'd4283090, -25'd1620629}}, '{'{25'd3009739, -25'd3974399, -25'd3897226, -25'd3704294, 25'd3511362, 25'd2893980, 25'd3241257, -25'd3048325, 25'd964660}, '{25'd3279844, -25'd501623, 25'd655969, -25'd424450, -25'd2392357, 25'd3279844, -25'd3897226, -25'd1659215, 25'd3549949}, '{25'd1697801, -25'd3318430, -25'd1041833, -25'd4012985, -25'd1620629, -25'd1852147, -25'd2816807, 25'd1003246, -25'd887487}, '{-25'd848901, -25'd3125498, -25'd2083665, 25'd4591781, 25'd3357017, -25'd463037, 25'd3665708, 25'd4090158, 25'd3357017}, '{25'd2816807, -25'd3048325, -25'd3820053, -25'd617382, -25'd1890733, 25'd2508116, 25'd3627121, 25'd1350524, -25'd2392357}, '{-25'd3742881, 25'd0, 25'd2585289, 25'd4244504, -25'd3627121, -25'd1543456, 25'd4476022, 25'd578796, -25'd2508116}, '{25'd4205917, 25'd3241257, -25'd3202671, -25'd2238011, 25'd2315184, -25'd1041833, 25'd2315184, -25'd3511362, 25'd2315184}, '{-25'd2083665, 25'd2546702, 25'd3665708, 25'd2778221, -25'd2353770, -25'd1311938, 25'd3549949, -25'd2430943, -25'd540210}, '{25'd2739634, 25'd4012985, -25'd1350524, -25'd270105, 25'd1080419, -25'd540210, -25'd2083665, 25'd1427697, 25'd1234765}}, '{'{-25'd2585289, -25'd2045079, -25'd1003246, 25'd3318430, 25'd3318430, -25'd1929320, -25'd3164085, 25'd4128745, -25'd2469529}, '{-25'd3704294, -25'd964660, -25'd2469529, 25'd4321677, 25'd0, 25'd2122252, 25'd1774974, -25'd3665708, -25'd4012985}, '{25'd1504870, -25'd4051572, -25'd3588535, 25'd1041833, -25'd2006493, 25'd1504870, -25'd2353770, 25'd1003246, -25'd192932}, '{25'd424450, -25'd2816807, 25'd4090158, 25'd1080419, 25'd4668954, 25'd2585289, -25'd3820053, -25'd1119006, 25'd270105}, '{-25'd1967906, -25'd77173, 25'd1929320, -25'd2546702, 25'd4900473, -25'd1659215, 25'd2739634, 25'd4668954, -25'd3781467}, '{-25'd1543456, 25'd2546702, -25'd2585289, -25'd2971153, -25'd1157592, 25'd347278, -25'd463037, -25'd2508116, 25'd192932}, '{25'd1659215, -25'd1697801, 25'd964660, 25'd1736388, 25'd694555, -25'd2315184, -25'd1080419, 25'd3742881, 25'd2199425}, '{-25'd578796, 25'd1852147, 25'd3318430, -25'd154346, 25'd3434189, 25'd4012985, 25'd2199425, -25'd1041833, -25'd2469529}, '{25'd887487, 25'd4321677, -25'd3935813, -25'd3974399, -25'd1350524, -25'd3897226, -25'd578796, 25'd1157592, -25'd1080419}}},
    '{'{'{-25'd1231128, -25'd2234270, 25'd3191814, 25'd3784579, 25'd2371062, 25'd364779, -25'd364779, 25'd3328606, 25'd1778296}, '{25'd3146217, 25'd0, 25'd1185531, 25'd4878916, 25'd775155, -25'd957544, 25'd1687102, -25'd1778296, -25'd1367920}, '{25'd273584, -25'd2143075, -25'd2918230, -25'd319181, 25'd2507854, -25'd1504712, 25'd2781438, 25'd4605331, -25'd3055022}, '{25'd820752, 25'd2553451, -25'd2507854, 25'd4878916, 25'd1139934, 25'd1732699, 25'd1276726, -25'd3283009, 25'd1459115}, '{-25'd1459115, -25'd227987, 25'd4650929, 25'd1231128, -25'd4058163, -25'd4696526, -25'd1960686, -25'd227987, -25'd319181}, '{25'd3146217, -25'd1367920, -25'd2188672, -25'd1504712, 25'd1413518, 25'd91195, -25'd3328606, 25'd3191814, -25'd3510995}, '{25'd4696526, 25'd3875774, -25'd2097478, -25'd3283009, 25'd2735840, -25'd866349, 25'd3556593, -25'd3647787, 25'd5152500}, '{25'd3283009, -25'd1641504, 25'd5061305, -25'd1413518, -25'd1778296, -25'd3465398, -25'd683960, 25'd3100619, 25'd2599048}, '{-25'd2918230, 25'd4103761, 25'd3556593, -25'd1094336, 25'd957544, 25'd4103761, 25'd957544, -25'd2188672, 25'd5243694}}, '{'{25'd5061305, -25'd2644646, -25'd227987, -25'd1595907, 25'd1276726, -25'd2599048, 25'd45597, 25'd1139934, 25'd1595907}, '{25'd2553451, 25'd3055022, 25'd3738982, -25'd1550310, -25'd2097478, 25'd3419801, -25'd182389, -25'd1094336, -25'd1778296}, '{-25'd1139934, 25'd4878916, 25'd4650929, -25'd2279867, -25'd2507854, -25'd1413518, -25'd683960, -25'd683960, -25'd1595907}, '{25'd5243694, -25'd364779, 25'd2827035, 25'd820752, 25'd4331747, -25'd4149358, 25'd2553451, -25'd1550310, -25'd957544}, '{-25'd2781438, 25'd3693385, 25'd364779, 25'd775155, -25'd3191814, -25'd1823894, -25'd1687102, 25'd638363, -25'd2827035}, '{25'd3510995, 25'd2690243, 25'd4377345, -25'd1915088, -25'd3693385, -25'd2599048, -25'd3055022, 25'd2599048, 25'd5015708}, '{25'd2553451, 25'd501571, -25'd638363, 25'd592765, -25'd1550310, 25'd273584, 25'd1641504, 25'd957544, -25'd182389}, '{25'd5790862, -25'd1732699, 25'd2963827, 25'd3693385, 25'd4012566, -25'd4012566, -25'd3009425, -25'd1550310, 25'd319181}, '{-25'd1960686, 25'd2553451, -25'd1732699, 25'd5152500, 25'd1276726, 25'd2234270, 25'd3191814, -25'd1915088, -25'd2872633}}, '{'{-25'd364779, 25'd866349, 25'd227987, 25'd911947, -25'd364779, 25'd2279867, -25'd3602190, -25'd3465398, -25'd729557}, '{-25'd3009425, 25'd4559734, 25'd911947, 25'd2279867, -25'd273584, 25'd3100619, 25'd2963827, -25'd729557, -25'd820752}, '{25'd2325464, 25'd5426084, -25'd410376, 25'd3921371, -25'd547168, -25'd364779, 25'd2462256, 25'd227987, -25'd866349}, '{25'd136792, 25'd3830177, 25'd5745265, 25'd1367920, 25'd2371062, -25'd1413518, 25'd45597, 25'd2553451, -25'd2507854}, '{-25'd775155, 25'd3374203, 25'd3921371, -25'd1550310, 25'd45597, -25'd1231128, -25'd4286150, 25'd4559734, 25'd4787721}, '{25'd592765, 25'd4924513, 25'd1915088, -25'd3647787, 25'd1276726, 25'd3146217, -25'd1869491, -25'd1550310, 25'd4559734}, '{-25'd547168, 25'd2918230, 25'd501571, -25'd2006283, 25'd2553451, -25'd2553451, 25'd45597, 25'd866349, 25'd364779}, '{25'd4787721, 25'd911947, 25'd2507854, 25'd957544, 25'd2051880, -25'd3784579, 25'd2918230, -25'd136792, -25'd1915088}, '{-25'd45597, 25'd5334889, 25'd729557, 25'd957544, 25'd683960, 25'd4787721, -25'd1231128, -25'd1778296, 25'd1778296}}},
    '{'{'{25'd1641007, 25'd2974325, -25'd3897392, -25'd717941, 25'd1264943, -25'd1367506, -25'd3452952, -25'd1128192, 25'd3179451}, '{-25'd615378, -25'd1094005, -25'd820503, 25'd1538444, 25'd2632449, 25'd2290572, 25'd3726453, 25'd3042700, -25'd136751}, '{25'd307689, 25'd3931579, -25'd1504256, 25'd2290572, -25'd1504256, 25'd1470069, -25'd957254, 25'd102563, -25'd1196568}, '{-25'd1059817, 25'd3008513, -25'd2529886, 25'd752128, 25'd2974325, -25'd2666636, 25'd3555515, 25'd1230755, -25'd273501}, '{25'd376064, 25'd2017071, 25'd3350389, 25'd410252, -25'd615378, 25'd2598261, -25'd1606819, -25'd1846133, 25'd1606819}, '{25'd1504256, -25'd3350389, -25'd1641007, 25'd1538444, 25'd2051259, -25'd3487140, 25'd3999954, -25'd2153822, 25'd2461510}, '{-25'd1914508, -25'd478627, 25'd3452952, -25'd1162380, -25'd478627, -25'd1401693, -25'd2837575, -25'd1162380, 25'd2051259}, '{-25'd786316, 25'd2188009, -25'd2393135, 25'd649565, 25'd4239268, 25'd820503, 25'd1538444, -25'd1811945, 25'd2871762}, '{25'd3726453, 25'd2632449, 25'd3897392, -25'd3863204, -25'd3350389, 25'd1059817, 25'd3794829, -25'd4239268, 25'd2358948}}, '{'{25'd2837575, 25'd3111076, 25'd2974325, -25'd239314, 25'd2188009, -25'd3213639, 25'd683753, 25'd1811945, -25'd2837575}, '{25'd307689, -25'd3247826, 25'd136751, -25'd581190, -25'd205126, -25'd1128192, 25'd3282014, -25'd2085446, -25'd1948696}, '{-25'd136751, -25'd3999954, 25'd2085446, -25'd2051259, 25'd2666636, -25'd205126, 25'd444439, -25'd1743570, -25'd683753}, '{-25'd341876, 25'd1914508, -25'd1675195, -25'd1504256, 25'd2119634, -25'd1059817, -25'd1299131, 25'd3555515, -25'd2256385}, '{25'd3213639, 25'd1059817, 25'd1094005, -25'd2632449, -25'd2461510, 25'd4341831, 25'd3179451, 25'd4341831, -25'd3589703}, '{25'd4239268, -25'd1504256, 25'd3316202, -25'd1675195, 25'd1914508, 25'd2940137, 25'd2461510, 25'd1504256, -25'd3316202}, '{25'd1914508, 25'd649565, 25'd3760641, -25'd1196568, 25'd3452952, -25'd1538444, -25'd1572632, -25'd2940137, 25'd1059817}, '{25'd4034142, 25'd3897392, 25'd1162380, 25'd2051259, 25'd1094005, 25'd341876, -25'd2495698, 25'd444439, 25'd444439}, '{25'd2598261, 25'd1264943, 25'd3965767, -25'd1538444, -25'd3487140, 25'd2598261, -25'd2017071, 25'd1196568, 25'd1606819}}, '{'{-25'd2358948, -25'd1538444, 25'd3897392, -25'd273501, 25'd4170893, 25'd547002, 25'd2598261, -25'd1025629, 25'd2085446}, '{-25'd136751, -25'd3384577, 25'd3145263, 25'd3829016, -25'd3418765, -25'd2119634, 25'd1299131, -25'd2290572, -25'd1948696}, '{-25'd991442, -25'd1880320, 25'd1504256, 25'd376064, -25'd1435881, 25'd3213639, 25'd4136705, -25'd2153822, 25'd1914508}, '{25'd1777758, 25'd2358948, -25'd3316202, 25'd1196568, 25'd1401693, -25'd4034142, -25'd4034142, 25'd3794829, -25'd68375}, '{-25'd1709382, -25'd1948696, 25'd1606819, -25'd2700824, -25'd786316, -25'd1128192, -25'd1094005, 25'd4273456, -25'd1777758}, '{-25'd3623890, -25'd3282014, 25'd1641007, -25'd3042700, 25'd752128, -25'd3179451, 25'd683753, 25'd2290572, 25'd683753}, '{25'd3521327, 25'd581190, -25'd3350389, 25'd957254, 25'd3316202, -25'd683753, 25'd1982883, 25'd2222197, 25'd3794829}, '{25'd923066, 25'd512815, 25'd3658078, -25'd1059817, -25'd478627, 25'd2153822, 25'd1948696, 25'd3384577, 25'd1675195}, '{-25'd136751, -25'd3931579, -25'd3999954, -25'd4068330, -25'd3316202, 25'd3418765, 25'd1333318, 25'd3623890, -25'd3692266}}},
    '{'{'{-25'd125540, 25'd2636339, 25'd0, -25'd8160095, -25'd753240, 25'd2761878, -25'd3515118, 25'd125540, -25'd1255399}, '{25'd2887418, 25'd753240, -25'd7532396, -25'd8411175, -25'd2761878, 25'd3264038, -25'd2887418, -25'd3640658, -25'd1506479}, '{-25'd1129859, -25'd4519437, -25'd5021597, -25'd7155776, 25'd1004319, 25'd2636339, 25'd1004319, -25'd376620, 25'd3389578}, '{-25'd7030236, -25'd6025917, 25'd1506479, 25'd1883099, 25'd9289955, 25'd1004319, -25'd2510799, 25'd502160, 25'd2134179}, '{-25'd6779156, -25'd2008639, 25'd1757559, 25'd2636339, 25'd15190332, 25'd8160095, 25'd3138498, -25'd376620, -25'd125540}, '{-25'd2134179, 25'd1632019, -25'd125540, 25'd1506479, 25'd15943571, 25'd4519437, 25'd5649297, -25'd251080, -25'd2259719}, '{-25'd3138498, -25'd5147137, 25'd753240, 25'd125540, 25'd13432773, 25'd9038875, 25'd4644977, -25'd3389578, -25'd878780}, '{-25'd1129859, -25'd3389578, -25'd3389578, 25'd2385259, 25'd3389578, 25'd5774837, -25'd1883099, -25'd1004319, 25'd1380939}, '{25'd753240, 25'd1632019, 25'd1506479, -25'd1129859, 25'd3640658, 25'd2134179, 25'd3138498, -25'd1004319, 25'd2761878}}, '{'{-25'd502160, -25'd1632019, -25'd6025917, -25'd4519437, 25'd3138498, -25'd1255399, -25'd1380939, 25'd2385259, 25'd3264038}, '{25'd4770517, -25'd2385259, -25'd2134179, -25'd8913335, 25'd5649297, -25'd1004319, 25'd3389578, 25'd4770517, 25'd6779156}, '{25'd3515118, 25'd376620, -25'd4770517, -25'd7657936, 25'd1632019, 25'd1129859, -25'd2008639, 25'd2761878, 25'd376620}, '{-25'd4393898, -25'd4017278, 25'd2887418, -25'd2761878, 25'd9164415, -25'd251080, -25'd5021597, -25'd753240, 25'd2134179}, '{-25'd4519437, -25'd4770517, 25'd4142818, 25'd4770517, 25'd10670894, 25'd7406856, 25'd2259719, -25'd1506479, 25'd627700}, '{-25'd3012958, -25'd4268358, 25'd5900377, 25'd6779156, 25'd11298594, 25'd4770517, -25'd5900377, -25'd4393898, -25'd5147137}, '{-25'd2761878, -25'd3012958, -25'd1129859, 25'd1883099, 25'd11549674, 25'd3138498, -25'd4896057, -25'd6402536, -25'd5398217}, '{-25'd251080, -25'd1757559, -25'd502160, 25'd1632019, 25'd125540, 25'd627700, -25'd4770517, -25'd5900377, -25'd1506479}, '{25'd3389578, -25'd1757559, -25'd1883099, -25'd3515118, 25'd1506479, 25'd1883099, 25'd0, -25'd627700, 25'd6151457}}, '{'{25'd6528076, 25'd3012958, -25'd125540, -25'd8913335, 25'd2636339, 25'd8536715, 25'd5147137, 25'd8034556, 25'd3640658}, '{25'd3766198, 25'd2385259, -25'd1757559, -25'd4896057, 25'd3012958, 25'd2385259, -25'd1129859, 25'd4896057, 25'd7783476}, '{25'd376620, -25'd4268358, -25'd4268358, -25'd9666575, 25'd2761878, -25'd3389578, -25'd125540, -25'd627700, 25'd1883099}, '{25'd878780, -25'd4519437, -25'd7281316, -25'd6653616, 25'd6653616, 25'd4142818, 25'd3012958, 25'd1757559, -25'd1506479}, '{-25'd1255399, -25'd5272677, -25'd3515118, -25'd1506479, 25'd7406856, 25'd4896057, -25'd2887418, -25'd4142818, -25'd753240}, '{-25'd4770517, 25'd0, 25'd2008639, 25'd1757559, 25'd14813712, 25'd8662255, 25'd5147137, -25'd4142818, -25'd1757559}, '{25'd0, -25'd1380939, -25'd3515118, 25'd4770517, 25'd8787795, 25'd1506479, -25'd4142818, 25'd1506479, -25'd2008639}, '{-25'd125540, -25'd6276997, 25'd125540, -25'd1632019, 25'd2510799, 25'd5900377, 25'd627700, -25'd2008639, -25'd251080}, '{-25'd753240, -25'd4017278, -25'd3138498, -25'd627700, -25'd1004319, -25'd3264038, -25'd4896057, 25'd2636339, 25'd5398217}}},
    '{'{'{25'd1774768, -25'd6263886, -25'd2714351, -25'd11066199, 25'd208796, 25'd4384720, -25'd2505555, -25'd1565972, -25'd313194}, '{-25'd2401156, -25'd10022218, -25'd13154161, -25'd11692588, 25'd1252777, -25'd5115507, -25'd2296758, -25'd5533100, -25'd3549536}, '{-25'd9500228, -25'd11796986, -25'd7203469, -25'd12110180, 25'd1461573, 25'd1983564, 25'd835185, -25'd313194, -25'd5533100}, '{-25'd10753005, -25'd13362958, -25'd7412266, -25'd2818749, 25'd3758332, 25'd313194, -25'd521991, -25'd3027545, -25'd8351848}, '{25'd2609953, 25'd3027545, 25'd5115507, 25'd6785877, 25'd9813422, 25'd8873839, 25'd9813422, 25'd1565972, 25'd1670370}, '{25'd2087962, 25'd8560645, 25'd3236341, 25'd3340739, 25'd11274995, 25'd2401156, 25'd1983564, 25'd5115507, 25'd6681479}, '{25'd4697915, 25'd3862730, 25'd208796, 25'd5428702, 25'd1670370, 25'd1252777, 25'd6368284, -25'd1357175, 25'd5846294}, '{25'd6055090, -25'd1148379, -25'd2714351, -25'd313194, 25'd4489119, 25'd1357175, -25'd730787, 25'd2609953, 25'd1774768}, '{25'd3862730, -25'd835185, -25'd4384720, 25'd2192360, 25'd104398, 25'd6055090, 25'd3236341, 25'd7307867, 25'd2087962}}, '{'{-25'd1461573, -25'd5219905, 25'd939583, -25'd6159488, 25'd3131943, 25'd104398, 25'd6159488, 25'd626389, 25'd4697915}, '{-25'd8247450, -25'd5741896, -25'd9709024, -25'd7516664, -25'd521991, 25'd3653934, 25'd730787, -25'd2192360, 25'd1148379}, '{-25'd5533100, -25'd8769441, -25'd7099071, -25'd2087962, -25'd1357175, 25'd4593517, -25'd626389, 25'd2609953, 25'd2192360}, '{-25'd10126616, -25'd5533100, -25'd10961801, -25'd5219905, -25'd1252777, -25'd730787, -25'd1983564, -25'd3653934, -25'd7099071}, '{25'd4071526, 25'd417592, 25'd5219905, 25'd1774768, 25'd8143052, 25'd7934256, 25'd2505555, 25'd7621062, 25'd1148379}, '{25'd3236341, 25'd1879166, 25'd2609953, 25'd0, 25'd10857403, 25'd1983564, 25'd4489119, 25'd2609953, 25'd2192360}, '{-25'd626389, -25'd1774768, 25'd2296758, -25'd417592, 25'd835185, -25'd1565972, 25'd730787, 25'd5011109, 25'd2609953}, '{-25'd2401156, 25'd1043981, -25'd313194, -25'd6785877, 25'd1774768, -25'd2296758, 25'd939583, -25'd2192360, 25'd835185}, '{25'd313194, -25'd6263886, -25'd1983564, -25'd1983564, 25'd2087962, -25'd3967128, -25'd208796, 25'd3967128, 25'd3131943}}, '{'{25'd5846294, -25'd2401156, -25'd1983564, -25'd4802313, 25'd104398, 25'd2296758, 25'd3236341, 25'd2714351, -25'd2087962}, '{-25'd1252777, -25'd4384720, -25'd8560645, -25'd3027545, -25'd4384720, 25'd2087962, 25'd1043981, -25'd3758332, -25'd835185}, '{-25'd5846294, -25'd4593517, -25'd8143052, -25'd4384720, -25'd1670370, 25'd1774768, -25'd6263886, -25'd1565972, 25'd0}, '{-25'd1357175, -25'd7829858, -25'd5533100, -25'd7203469, -25'd1252777, 25'd208796, -25'd1983564, -25'd5950692, -25'd6577081}, '{25'd7516664, 25'd4802313, 25'd7099071, 25'd2296758, 25'd7412266, 25'd3549536, 25'd6368284, 25'd2818749, -25'd208796}, '{25'd2192360, 25'd8351848, 25'd7203469, 25'd521991, 25'd7934256, 25'd2087962, 25'd4802313, 25'd3445138, -25'd1565972}, '{25'd6890275, 25'd5950692, 25'd5428702, 25'd5011109, 25'd5846294, 25'd4071526, -25'd1983564, -25'd2401156, 25'd208796}, '{25'd1670370, 25'd5115507, -25'd1252777, -25'd3027545, 25'd3340739, -25'd3653934, 25'd1565972, 25'd3236341, -25'd3340739}, '{25'd3758332, 25'd2087962, 25'd1670370, -25'd7307867, 25'd1565972, 25'd939583, -25'd5115507, 25'd2714351, 25'd4071526}}},
    '{'{'{-25'd1074447, 25'd3509861, -25'd3939640, 25'd3760565, -25'd1934005, 25'd859558, 25'd4226159, 25'd2793563, 25'd2865192}, '{25'd2686118, -25'd1683301, 25'd1110262, 25'd1432596, 25'd322334, 25'd4441048, -25'd2614488, -25'd3868010, 25'd0}, '{-25'd1253522, 25'd1719115, -25'd358149, -25'd1575856, -25'd2113079, -25'd107445, -25'd3044267, -25'd1360966, 25'd2363784}, '{-25'd608853, 25'd3402416, -25'd967002, 25'd1898190, -25'd3330786, 25'd2721933, 25'd1217707, 25'd2829378, 25'd787928}, '{-25'd501409, 25'd1396781, 25'd1826560, -25'd2793563, 25'd2005635, 25'd4226159, 25'd1504226, -25'd2901007, -25'd2148894}, '{25'd3115897, 25'd322334, -25'd1325152, 25'd752113, 25'd1504226, 25'd716298, 25'd1969820, 25'd3903825, -25'd3187527}, '{-25'd644668, -25'd465594, 25'd2041450, -25'd3080082, 25'd4261974, -25'd895373, -25'd1540041, -25'd3724750, -25'd3008452}, '{25'd4441048, 25'd4190344, -25'd716298, -25'd2041450, -25'd680483, 25'd1002817, 25'd2113079, -25'd608853, 25'd2220524}, '{-25'd286519, 25'd1611671, -25'd1969820, -25'd1360966, -25'd2650303, -25'd2578673, -25'd2829378, -25'd2721933, 25'd3975455}}, '{'{25'd393964, -25'd250704, -25'd573038, 25'd322334, -25'd3653120, -25'd35815, 25'd3868010, 25'd4082899, -25'd1504226}, '{-25'd2507043, 25'd429779, 25'd2327969, -25'd3402416, -25'd3008452, -25'd1969820, -25'd1253522, -25'd3438231, 25'd823743}, '{-25'd1002817, -25'd35815, -25'd2686118, -25'd1038632, 25'd1826560, 25'd859558, -25'd2471229, 25'd1217707, 25'd2721933}, '{25'd4441048, -25'd179075, -25'd1934005, 25'd2686118, 25'd1468411, -25'd71630, -25'd2757748, 25'd3438231, -25'd1074447}, '{-25'd250704, 25'd2901007, -25'd107445, 25'd2972637, -25'd1862375, -25'd3187527, -25'd2077265, -25'd3187527, -25'd2793563}, '{25'd3259156, 25'd4011269, -25'd2399599, -25'd2793563, -25'd716298, 25'd3115897, 25'd3796380, 25'd3223342, 25'd967002}, '{25'd3760565, -25'd214889, -25'd358149, 25'd1826560, 25'd1790745, 25'd1504226, -25'd3115897, 25'd2363784, 25'd2113079}, '{-25'd3115897, 25'd2578673, 25'd2292154, -25'd3438231, 25'd2542858, -25'd71630, -25'd787928, -25'd787928, 25'd4333604}, '{-25'd1432596, 25'd4548493, 25'd1146077, -25'd3796380, -25'd429779, -25'd3115897, 25'd4226159, -25'd1540041, -25'd3044267}}, '{'{-25'd2542858, 25'd4154529, -25'd1038632, -25'd1719115, -25'd1038632, 25'd2901007, 25'd3688935, -25'd1575856, 25'd2578673}, '{-25'd1754930, -25'd1719115, 25'd4226159, 25'd107445, -25'd1754930, 25'd859558, 25'd179075, -25'd1934005, 25'd286519}, '{25'd2363784, 25'd823743, 25'd1611671, -25'd3402416, 25'd3545676, 25'd1862375, -25'd2972637, -25'd322334, 25'd1575856}, '{25'd3044267, 25'd2005635, 25'd3939640, 25'd322334, 25'd250704, 25'd1754930, 25'd1110262, 25'd1074447, 25'd2220524}, '{-25'd3223342, 25'd2901007, 25'd4154529, -25'd2578673, 25'd1719115, 25'd1468411, -25'd3760565, 25'd4512678, -25'd3509861}, '{25'd4441048, -25'd1002817, -25'd3080082, 25'd1038632, 25'd895373, 25'd859558, -25'd3474046, -25'd1790745, -25'd1575856}, '{25'd214889, 25'd3903825, -25'd1969820, 25'd2757748, 25'd2399599, 25'd3939640, 25'd3653120, -25'd1898190, -25'd2327969}, '{-25'd859558, 25'd2005635, 25'd3223342, -25'd2363784, -25'd2184709, -25'd3080082, -25'd716298, 25'd1862375, -25'd2292154}, '{25'd3975455, 25'd1611671, -25'd1253522, 25'd4512678, 25'd179075, -25'd1360966, 25'd3294971, -25'd2614488, 25'd752113}}},
    '{'{'{-25'd3612723, 25'd4452043, -25'd2226021, -25'd328429, 25'd3612723, 25'd2408482, -25'd3649215, -25'd3357278, -25'd547382}, '{25'd3211309, -25'd1350210, -25'd693351, -25'd583874, -25'd2809896, -25'd3904660, 25'd2335498, -25'd839319, -25'd2371990}, '{25'd839319, -25'd3795184, 25'd1350210, -25'd36492, -25'd693351, 25'd0, 25'd4488535, 25'd4342566, -25'd3393770}, '{25'd3466754, -25'd1277225, -25'd364922, -25'd3722200, 25'd1240733, -25'd2408482, -25'd1496178, 25'd328429, -25'd2444974}, '{-25'd510890, -25'd766335, -25'd1861100, -25'd3612723, 25'd3539739, -25'd875812, 25'd2919372, -25'd3174817, 25'd620367}, '{-25'd3977645, -25'd2043561, 25'd1131257, -25'd839319, -25'd766335, 25'd2663927, 25'd2590943, 25'd4160105, -25'd2773404}, '{25'd1058272, -25'd3028849, -25'd1751623, 25'd547382, 25'd4233090, -25'd510890, 25'd109476, -25'd3941152, -25'd1423194}, '{-25'd839319, 25'd1788115, 25'd3977645, 25'd4050629, 25'd1824608, 25'd2153037, 25'd182461, 25'd583874, 25'd3357278}, '{25'd3284294, 25'd2700419, 25'd3685707, 25'd437906, 25'd3977645, -25'd3722200, 25'd3247802, -25'd1569163, 25'd1970576}}, '{'{-25'd1532670, 25'd2299006, 25'd437906, 25'd3284294, 25'd875812, -25'd1605655, -25'd3831676, 25'd1678639, 25'd3101833}, '{-25'd3649215, 25'd2335498, 25'd3685707, -25'd1715131, 25'd328429, 25'd2262513, 25'd1277225, -25'd1021780, -25'd2554451}, '{25'd4160105, 25'd2846388, 25'd2627435, -25'd2481466, 25'd3101833, 25'd3868168, 25'd4415550, 25'd218953, -25'd437906}, '{-25'd3174817, -25'd1240733, 25'd328429, -25'd291937, -25'd839319, 25'd802827, 25'd36492, -25'd1204241, -25'd839319}, '{-25'd1715131, -25'd839319, -25'd364922, 25'd3320786, 25'd2590943, 25'd3284294, -25'd3138325, -25'd36492, -25'd3211309}, '{25'd2007068, 25'd3539739, 25'd3393770, 25'd1861100, -25'd2700419, 25'd1240733, 25'd1788115, -25'd3284294, -25'd1897592}, '{-25'd3430262, -25'd583874, -25'd2919372, -25'd3831676, -25'd2554451, 25'd3868168, -25'd3612723, -25'd729843, 25'd1532670}, '{-25'd1313717, -25'd4123613, 25'd3977645, -25'd3138325, 25'd2773404, -25'd1605655, 25'd2882880, -25'd2299006, -25'd2262513}, '{-25'd182461, 25'd1934084, 25'd3868168, 25'd1277225, -25'd255445, 25'd656859, -25'd547382, 25'd1313717, 25'd3904660}}, '{'{-25'd1386702, -25'd145969, 25'd4634503, -25'd2992356, 25'd36492, -25'd2992356, 25'd2554451, -25'd1423194, 25'd2517958}, '{25'd4087121, 25'd1897592, 25'd4160105, -25'd2153037, 25'd802827, 25'd4415550, -25'd1021780, 25'd1569163, 25'd255445}, '{25'd4634503, 25'd1094765, 25'd3138325, 25'd474398, 25'd2481466, -25'd1605655, 25'd3539739, -25'd2371990, -25'd1715131}, '{-25'd36492, -25'd3539739, -25'd1167749, -25'd3758692, -25'd2809896, 25'd4598011, 25'd766335, -25'd620367, -25'd1021780}, '{25'd3211309, 25'd620367, 25'd3649215, 25'd3065341, 25'd2262513, -25'd1788115, 25'd1459686, -25'd2153037, 25'd3503247}, '{-25'd1058272, 25'd2371990, 25'd2262513, 25'd2846388, 25'd4488535, 25'd1386702, 25'd2080053, -25'd2846388, -25'd2043561}, '{-25'd766335, 25'd1094765, -25'd1642147, -25'd2846388, -25'd2846388, -25'd1605655, 25'd1751623, 25'd3211309, -25'd3393770}, '{25'd4087121, 25'd4014137, 25'd1532670, -25'd620367, 25'd1751623, 25'd1824608, 25'd2919372, -25'd1751623, 25'd4050629}, '{-25'd2226021, 25'd4525027, -25'd291937, 25'd2408482, 25'd2043561, 25'd3868168, 25'd4379058, -25'd328429, 25'd2408482}}},
    '{'{'{25'd3149477, 25'd1861054, -25'd2505266, -25'd3614740, -25'd572632, 25'd1574738, -25'd1717896, -25'd1932633, 25'd2075791}, '{25'd3364214, 25'd4187372, 25'd1968423, -25'd1252633, -25'd178948, 25'd2648424, 25'd536843, 25'd3006319, -25'd1861054}, '{25'd1181054, -25'd1538949, 25'd930527, -25'd1324212, -25'd4151583, -25'd4115793, 25'd3400003, 25'd1109475, 25'd1538949}, '{-25'd143158, -25'd2755792, 25'd1896844, -25'd3901056, 25'd823159, 25'd3507372, 25'd3077898, 25'd2397897, 25'd71579}, '{25'd536843, 25'd3865267, -25'd2326318, -25'd1717896, -25'd1431580, 25'd2075791, 25'd2290529, 25'd2147371, -25'd2970529}, '{25'd894738, 25'd3972635, 25'd4223162, -25'd3328424, 25'd3328424, -25'd2004212, -25'd3614740, -25'd501053, -25'd3006319}, '{-25'd3292635, 25'd644211, -25'd3865267, 25'd1503159, 25'd1288422, 25'd2612634, -25'd715790, -25'd1682107, 25'd1109475}, '{25'd2827371, -25'd322106, 25'd1574738, 25'd1610528, 25'd1288422, -25'd4151583, 25'd1431580, -25'd286316, -25'd3400003}, '{-25'd2362108, -25'd572632, -25'd2612634, 25'd250527, -25'd1932633, 25'd4115793, -25'd2183160, 25'd3364214, 25'd322106}}, '{'{25'd4545268, 25'd3042108, 25'd107369, -25'd3113687, 25'd1968423, -25'd2648424, 25'd286316, 25'd0, 25'd4437899}, '{-25'd1181054, -25'd3507372, 25'd4258951, 25'd1109475, -25'd2684213, 25'd2827371, 25'd143158, 25'd715790, -25'd3185266}, '{25'd4473689, -25'd3543161, 25'd1538949, -25'd3292635, 25'd3256845, 25'd3543161, 25'd250527, -25'd3578951, -25'd2791582}, '{-25'd2469476, -25'd1288422, -25'd1610528, 25'd3865267, 25'd107369, -25'd894738, -25'd3901056, 25'd4080004, -25'd2290529}, '{25'd823159, 25'd3364214, 25'd2541055, 25'd894738, -25'd1932633, -25'd501053, -25'd1216843, -25'd2612634, -25'd787369}, '{25'd2469476, -25'd1431580, -25'd536843, 25'd930527, -25'd3793688, 25'd1073685, 25'd2111581, -25'd250527, 25'd4044214}, '{-25'd2075791, 25'd3972635, -25'd2183160, 25'd787369, -25'd715790, -25'd2183160, -25'd357895, -25'd1682107, 25'd322106}, '{-25'd322106, 25'd2648424, 25'd930527, -25'd2505266, 25'd1037896, -25'd1682107, 25'd1753686, 25'd1431580, -25'd2254739}, '{25'd4366320, 25'd3435793, 25'd3650530, -25'd3185266, -25'd1288422, -25'd1610528, 25'd3865267, 25'd536843, 25'd930527}}, '{'{25'd3077898, 25'd787369, -25'd2326318, -25'd1610528, -25'd2505266, 25'd4258951, -25'd4151583, 25'd286316, 25'd3829477}, '{25'd894738, 25'd4151583, 25'd393685, -25'd357895, 25'd2684213, -25'd1252633, -25'd3650530, 25'd1896844, 25'd680001}, '{25'd3936846, 25'd3578951, 25'd2254739, -25'd3185266, 25'd1646317, -25'd3113687, 25'd2254739, 25'd1073685, -25'd4044214}, '{25'd3328424, 25'd3865267, 25'd1610528, 25'd1252633, 25'd3113687, 25'd1431580, -25'd2326318, -25'd393685, -25'd357895}, '{-25'd1610528, 25'd3400003, 25'd1073685, -25'd3185266, 25'd1431580, -25'd1145264, -25'd3471582, 25'd1968423, 25'd1789475}, '{-25'd1538949, 25'd1288422, -25'd393685, -25'd1610528, 25'd4115793, -25'd3614740, 25'd1360001, 25'd787369, 25'd1538949}, '{-25'd1610528, 25'd1073685, -25'd1646317, -25'd3077898, 25'd1109475, 25'd465264, 25'd322106, -25'd966317, 25'd2004212}, '{-25'd357895, 25'd1216843, 25'd715790, 25'd3221056, -25'd2147371, 25'd751580, -25'd2254739, -25'd1216843, -25'd823159}, '{25'd1717896, -25'd2290529, -25'd3042108, -25'd3328424, 25'd4509478, 25'd1861054, -25'd2505266, -25'd3256845, 25'd4080004}}},
    '{'{'{25'd880592, -25'd3830575, 25'd4314901, 25'd4226841, 25'd3962664, -25'd1056710, -25'd3390279, 25'd3478338, 25'd3346249}, '{25'd220148, 25'd1717154, 25'd4050723, 25'd2333569, 25'd1276858, -25'd220148, 25'd132089, 25'd2157450, -25'd1232829}, '{-25'd1012681, 25'd1188799, -25'd132089, -25'd1585066, 25'd4446989, 25'd4446989, -25'd616414, 25'd2289539, 25'd1629095}, '{-25'd3214161, -25'd2861924, 25'd4667137, 25'd4270871, 25'd5195493, -25'd2245510, 25'd1937302, -25'd1012681, -25'd1717154}, '{-25'd1144770, -25'd2553717, 25'd3126101, -25'd528355, -25'd132089, -25'd396266, -25'd2597746, 25'd44030, 25'd3434309}, '{25'd1012681, -25'd2025362, 25'd0, 25'd1012681, 25'd1893273, -25'd308207, -25'd88059, 25'd704474, -25'd616414}, '{25'd2553717, 25'd4270871, 25'd3170131, 25'd1056710, -25'd1629095, -25'd1144770, 25'd3390279, 25'd3170131, 25'd1981332}, '{25'd220148, -25'd2333569, -25'd3126101, 25'd4623108, 25'd1541036, -25'd1893273, -25'd836562, -25'd176118, 25'd44030}, '{-25'd2289539, -25'd1761184, -25'd1144770, -25'd1761184, -25'd44030, -25'd1188799, 25'd1585066, -25'd4226841, 25'd572385}}, '{'{-25'd264178, -25'd3346249, 25'd3830575, -25'd1232829, 25'd2421628, -25'd4446989, 25'd3390279, 25'd176118, -25'd3478338}, '{-25'd3786545, 25'd2641776, 25'd528355, -25'd2465657, 25'd2113421, 25'd2025362, -25'd3038042, -25'd2817894, 25'd484326}, '{-25'd2157450, -25'd1981332, 25'd1012681, 25'd968651, -25'd1673125, 25'd1629095, 25'd2113421, 25'd2157450, 25'd2421628}, '{-25'd2861924, 25'd2641776, 25'd4270871, 25'd1276858, 25'd352237, -25'd2949983, -25'd1805214, 25'd1100740, -25'd2994013}, '{25'd528355, -25'd3610427, -25'd2685805, 25'd4006693, 25'd3214161, -25'd2465657, 25'd3258190, 25'd484326, -25'd1849243}, '{-25'd5063404, -25'd1408947, 25'd3566397, 25'd4623108, 25'd1188799, -25'd3698486, -25'd2905953, -25'd4182812, -25'd3786545}, '{-25'd4623108, 25'd1673125, -25'd2817894, -25'd2994013, -25'd1452977, 25'd1188799, 25'd2553717, -25'd3390279, 25'd352237}, '{25'd2861924, 25'd1232829, -25'd4711167, -25'd2025362, 25'd528355, 25'd2113421, -25'd1937302, 25'd1056710, 25'd1893273}, '{25'd924622, -25'd4402960, -25'd5063404, 25'd2994013, 25'd2553717, -25'd2025362, -25'd1056710, -25'd2994013, -25'd4887285}}, '{'{25'd2641776, -25'd1056710, 25'd1364918, -25'd2861924, 25'd2861924, -25'd1541036, 25'd3874605, 25'd1497006, 25'd3214161}, '{-25'd176118, -25'd748503, 25'd924622, -25'd660444, 25'd2773865, -25'd44030, 25'd3742516, 25'd4535049, 25'd1541036}, '{25'd396266, 25'd3654457, 25'd3346249, 25'd1364918, 25'd5151463, -25'd1673125, -25'd3170131, -25'd1717154, 25'd3786545}, '{25'd3214161, -25'd924622, -25'd396266, 25'd5591759, 25'd1144770, 25'd3610427, -25'd880592, -25'd2377598, 25'd44030}, '{-25'd1100740, 25'd5415641, 25'd1012681, 25'd5019374, 25'd3214161, 25'd5371611, 25'd2861924, -25'd704474, 25'd4887285}, '{25'd4535049, -25'd2333569, -25'd2157450, 25'd308207, 25'd2553717, 25'd3346249, 25'd3522368, 25'd3038042, 25'd880592}, '{25'd1849243, 25'd1144770, -25'd1056710, 25'd4138782, 25'd176118, 25'd220148, 25'd308207, 25'd1408947, -25'd2333569}, '{-25'd3962664, -25'd3918634, 25'd3478338, -25'd2377598, -25'd924622, -25'd1188799, 25'd352237, -25'd3698486, 25'd2069391}, '{25'd352237, -25'd704474, -25'd2157450, -25'd3302220, -25'd1276858, -25'd3390279, -25'd484326, -25'd1144770, 25'd2421628}}},
    '{'{'{-25'd3199452, 25'd186015, 25'd3943511, -25'd930073, -25'd446435, -25'd2827423, 25'd2157770, -25'd483638, -25'd3497076}, '{-25'd669653, 25'd4017917, -25'd1227697, -25'd2678611, 25'd3980714, 25'd2380988, -25'd1041682, 25'd2641408, -25'd2418191}, '{25'd1711335, 25'd1376509, -25'd260421, 25'd558044, -25'd297623, -25'd1302103, 25'd3869105, 25'd1860147, -25'd3236655}, '{-25'd1153291, 25'd1562523, -25'd1562523, 25'd2715814, 25'd595247, 25'd3087844, 25'd1078885, -25'd1450914, 25'd2641408}, '{-25'd2678611, 25'd3087844, 25'd334826, -25'd4166729, 25'd3199452, 25'd2827423, 25'd558044, -25'd372029, -25'd3236655}, '{25'd2008958, 25'd1153291, -25'd3385467, -25'd4501555, 25'd706856, -25'd1748538, -25'd297623, 25'd3608685, 25'd483638}, '{-25'd3720293, -25'd4092323, -25'd1711335, -25'd4278338, 25'd3311061, 25'd37203, 25'd1934553, 25'd1450914, -25'd2678611}, '{25'd3125047, 25'd297623, 25'd3683091, -25'd372029, -25'd2641408, -25'd3608685, -25'd1525320, 25'd1302103, 25'd520841}, '{-25'd111609, 25'd2976235, -25'd2083364, 25'd1860147, 25'd4055120, 25'd4092323, 25'd1748538, 25'd3013438, 25'd2083364}}, '{'{25'd2678611, 25'd3162249, 25'd2380988, -25'd3831902, 25'd2976235, -25'd2567003, 25'd2678611, 25'd781262, -25'd3273858}, '{25'd2418191, 25'd372029, -25'd4055120, 25'd3125047, -25'd744059, -25'd3311061, -25'd3534279, -25'd2939032, 25'd3720293}, '{-25'd3013438, -25'd4761976, 25'd1897350, -25'd483638, -25'd4538758, -25'd2790220, -25'd2083364, 25'd3906308, -25'd520841}, '{-25'd3645888, -25'd855668, 25'd2083364, 25'd3683091, -25'd2567003, 25'd1116088, 25'd74406, 25'd483638, -25'd3125047}, '{25'd1302103, -25'd4650367, -25'd2939032, -25'd2827423, 25'd2120567, -25'd2529800, 25'd3348264, -25'd1525320, -25'd3125047}, '{-25'd1116088, 25'd334826, 25'd1636929, 25'd1934553, 25'd1599726, -25'd74406, -25'd558044, -25'd2715814, 25'd3348264}, '{25'd2753017, 25'd2864626, -25'd3013438, 25'd223218, -25'd967276, 25'd1748538, 25'd520841, -25'd4017917, -25'd3125047}, '{-25'd4241135, -25'd1004479, 25'd3311061, -25'd669653, -25'd3273858, -25'd74406, -25'd3720293, 25'd2343785, -25'd74406}, '{-25'd3831902, -25'd2901829, -25'd3125047, -25'd3348264, -25'd3050641, -25'd260421, 25'd2380988, -25'd781262, 25'd3794699}}, '{'{25'd3348264, -25'd2269379, -25'd1302103, -25'd4538758, -25'd1860147, 25'd632450, 25'd2604205, 25'd148812, -25'd3497076}, '{25'd3348264, -25'd930073, 25'd2120567, -25'd2715814, -25'd2567003, -25'd669653, 25'd3199452, -25'd3348264, 25'd3459873}, '{-25'd4352743, 25'd744059, -25'd2641408, -25'd892870, 25'd223218, -25'd446435, 25'd1413712, -25'd2046161, 25'd446435}, '{25'd3236655, 25'd3348264, -25'd3125047, -25'd3013438, 25'd930073, 25'd3534279, -25'd2901829, 25'd1674132, 25'd3869105}, '{25'd297623, 25'd1376509, -25'd2083364, 25'd1525320, 25'd2641408, -25'd2678611, 25'd3087844, -25'd2120567, 25'd2343785}, '{-25'd930073, 25'd1153291, -25'd967276, -25'd4092323, -25'd4538758, -25'd1971756, 25'd1860147, -25'd4203932, -25'd706856}, '{25'd1822944, -25'd4129526, -25'd781262, 25'd3683091, -25'd3348264, -25'd3608685, -25'd4427149, -25'd1674132, -25'd2790220}, '{25'd2120567, -25'd744059, 25'd1934553, 25'd3683091, -25'd632450, 25'd3683091, -25'd37203, 25'd2455394, -25'd3459873}, '{25'd3645888, -25'd818465, -25'd3199452, 25'd3348264, -25'd632450, 25'd930073, 25'd4017917, 25'd2157770, -25'd2492597}}},
    '{'{'{-25'd1858765, 25'd3420127, -25'd3122725, 25'd3308601, -25'd3085550, -25'd817857, 25'd2713797, -25'd2974024, 25'd4200808}, '{25'd1524187, 25'd1561362, 25'd706331, 25'd2044641, -25'd1933115, -25'd3085550, 25'd2936848, -25'd3122725, 25'd1635713}, '{-25'd1784414, -25'd3643179, 25'd2565095, -25'd1895940, 25'd966558, -25'd966558, -25'd1561362, 25'd1672888, 25'd3568828}, '{-25'd1561362, -25'd1524187, 25'd2007466, 25'd2899673, 25'd4349510, -25'd1412661, -25'd2899673, 25'd2936848, 25'd1672888}, '{25'd2230518, 25'd2267693, 25'd3085550, 25'd520454, -25'd3606004, 25'd3271426, 25'd2899673, 25'd3680354, 25'd892207}, '{-25'd706331, -25'd1487012, 25'd1524187, 25'd4052107, 25'd2416394, 25'd2416394, -25'd1970291, 25'd2788147, -25'd1672888}, '{-25'd2304868, -25'd1412661, 25'd74351, -25'd3011199, -25'd2304868, 25'd669155, -25'd1858765, -25'd1412661, 25'd37175}, '{-25'd520454, -25'd3680354, 25'd557629, -25'd4423860, -25'd4609737, -25'd4386685, -25'd4758438, -25'd1858765, 25'd2193342}, '{25'd446104, -25'd260227, 25'd185876, 25'd706331, -25'd2118992, 25'd3085550, 25'd185876, -25'd966558, -25'd4014932}}, '{'{-25'd1710064, -25'd1635713, 25'd1895940, -25'd408928, 25'd3791880, -25'd37175, -25'd3420127, 25'd966558, 25'd3420127}, '{25'd2936848, 25'd4052107, 25'd1487012, 25'd3568828, -25'd4089283, 25'd1040908, 25'd74351, -25'd520454, -25'd1672888}, '{25'd1152434, -25'd892207, -25'd1895940, 25'd3606004, -25'd4163633, 25'd483279, 25'd4052107, -25'd520454, 25'd3568828}, '{25'd2490745, -25'd3494478, -25'd1895940, 25'd1635713, -25'd223052, -25'd2527920, 25'd4163633, 25'd3048374, 25'd1970291}, '{25'd817857, -25'd3717530, -25'd2193342, 25'd3345777, -25'd3643179, -25'd2825322, -25'd2342044, 25'd483279, -25'd483279}, '{-25'd2342044, 25'd966558, -25'd2342044, 25'd3940581, -25'd1301135, 25'd1970291, -25'd1933115, 25'd3940581, -25'd3866231}, '{25'd4349510, 25'd111526, 25'd706331, 25'd0, 25'd1672888, 25'd1672888, 25'd223052, -25'd2825322, 25'd2527920}, '{-25'd1858765, -25'd3717530, -25'd4237984, -25'd4721263, -25'd1412661, 25'd1635713, 25'd1449837, -25'd148701, -25'd483279}, '{25'd2342044, 25'd37175, -25'd111526, -25'd483279, -25'd2565095, 25'd37175, -25'd3606004, -25'd3606004, -25'd1263960}}, '{'{25'd2044641, 25'd4312334, -25'd297402, 25'd3643179, -25'd3829055, 25'd3680354, 25'd631980, -25'd3903406, 25'd297402}, '{-25'd483279, -25'd780681, -25'd3568828, -25'd2379219, -25'd1003733, -25'd3791880, 25'd483279, -25'd2304868, -25'd260227}, '{25'd2788147, -25'd260227, 25'd2118992, -25'd4498211, 25'd929382, 25'd4052107, 25'd1747239, -25'd3122725, -25'd1933115}, '{25'd223052, -25'd4163633, -25'd2974024, -25'd2862498, -25'd74351, 25'd2490745, 25'd1338311, 25'd1189609, -25'd892207}, '{25'd3680354, -25'd3308601, -25'd3717530, 25'd1672888, 25'd334578, -25'd1152434, -25'd706331, -25'd780681, -25'd3085550}, '{-25'd408928, -25'd4498211, -25'd855032, 25'd3085550, -25'd3159900, 25'd2118992, 25'd855032, -25'd1301135, -25'd2156167}, '{-25'd1933115, 25'd111526, -25'd1449837, 25'd260227, -25'd1821589, 25'd3011199, 25'd1487012, 25'd4126458, 25'd4535386}, '{25'd1226785, 25'd3048374, -25'd3308601, 25'd3717530, -25'd297402, 25'd2565095, 25'd37175, 25'd1933115, -25'd817857}, '{-25'd3606004, -25'd1635713, -25'd4014932, 25'd2007466, -25'd1933115, -25'd4052107, -25'd1858765, 25'd2342044, 25'd4349510}}},
    '{'{'{-25'd3539246, -25'd1408475, 25'd3719819, 25'd3972623, 25'd1950197, -25'd216689, -25'd3719819, -25'd469492, -25'd722295}, '{25'd1480705, 25'd2239115, 25'd3683705, 25'd2925295, 25'd2239115, -25'd505607, -25'd3358672, 25'd4044852, 25'd1841852}, '{-25'd2672492, -25'd2491918, 25'd3792049, -25'd1227902, -25'd613951, -25'd3467016, -25'd3214213, 25'd1047328, 25'd4514344}, '{-25'd1625164, -25'd1191787, 25'd3069754, 25'd3503131, -25'd1408475, -25'd1227902, 25'd3864278, 25'd794525, -25'd361148}, '{-25'd2383574, -25'd3900393, -25'd3322557, 25'd4044852, -25'd2203000, 25'd2058541, -25'd2997524, -25'd2203000, 25'd3178098}, '{25'd4080967, 25'd1877967, 25'd1300131, 25'd1769623, -25'd3430901, 25'd2961410, 25'd1877967, -25'd722295, 25'd3755934}, '{-25'd2708606, -25'd2311344, -25'd2816951, 25'd433377, 25'd541721, 25'd3214213, 25'd2455803, -25'd3972623, -25'd2058541}, '{25'd4333770, 25'd4333770, -25'd1372361, 25'd3322557, 25'd1155672, 25'd1661279, 25'd2708606, 25'd4044852, 25'd3033639}, '{-25'd3430901, 25'd0, 25'd2419688, -25'd2997524, 25'd3467016, -25'd361148, 25'd3033639, 25'd1841852, -25'd1733508}}, '{'{-25'd2419688, 25'd4442114, 25'd4514344, 25'd4153196, 25'd4406000, 25'd650066, -25'd3250328, -25'd2961410, 25'd613951}, '{25'd2203000, 25'd650066, -25'd3141983, -25'd2058541, 25'd1444590, 25'd2058541, -25'd2672492, -25'd3828164, 25'd3539246}, '{25'd1552934, 25'd2347459, -25'd2203000, 25'd4297655, 25'd1227902, 25'd2600262, 25'd4225426, 25'd4478229, -25'd2961410}, '{25'd469492, 25'd3105869, 25'd2058541, -25'd1408475, 25'd361148, -25'd252803, 25'd2997524, -25'd2997524, -25'd3683705}, '{-25'd938984, -25'd4044852, 25'd4261541, -25'd2744721, -25'd3755934, -25'd1697393, 25'd613951, 25'd4297655, -25'd2564147}, '{25'd686180, -25'd1047328, 25'd2780836, 25'd2130770, 25'd3467016, 25'd3105869, -25'd2022426, 25'd3033639, 25'd866754}, '{25'd2094656, 25'd1697393, 25'd3936508, -25'd3864278, -25'd3394787, 25'd3250328, 25'd1300131, 25'd3972623, -25'd3900393}, '{-25'd3322557, 25'd0, -25'd1661279, 25'd3503131, 25'd1914082, -25'd3828164, -25'd3214213, -25'd1914082, -25'd577836}, '{-25'd2419688, 25'd3105869, 25'd2311344, 25'd1914082, -25'd2889180, -25'd2744721, 25'd2889180, -25'd1047328, 25'd2853065}}, '{'{-25'd361148, 25'd3647590, -25'd2961410, 25'd830639, 25'd1516820, -25'd3430901, -25'd541721, -25'd3792049, -25'd722295}, '{25'd2347459, -25'd2961410, 25'd3539246, -25'd1372361, 25'd2961410, 25'd938984, -25'd1589049, 25'd2022426, 25'd2022426}, '{25'd1625164, -25'd3394787, 25'd4189311, -25'd3250328, -25'd3358672, 25'd1480705, -25'd1697393, 25'd0, 25'd2347459}, '{25'd3900393, -25'd794525, 25'd3178098, 25'd3141983, 25'd4514344, 25'd2130770, -25'd1155672, -25'd1408475, -25'd3864278}, '{25'd1372361, 25'd2311344, 25'd2636377, -25'd2130770, -25'd1805738, -25'd2780836, 25'd1011213, 25'd1372361, -25'd252803}, '{-25'd3683705, 25'd469492, -25'd2094656, 25'd3033639, 25'd4586573, 25'd2203000, -25'd3286442, -25'd2094656, 25'd2022426}, '{25'd2708606, -25'd1516820, 25'd2564147, -25'd1336246, -25'd1697393, -25'd3286442, 25'd3105869, -25'd686180, 25'd3394787}, '{-25'd433377, 25'd4080967, 25'd2311344, 25'd650066, 25'd397262, -25'd2419688, 25'd2780836, 25'd3394787, 25'd4297655}, '{25'd1372361, 25'd3864278, 25'd3611475, -25'd2600262, 25'd2744721, 25'd2239115, 25'd2455803, -25'd541721, -25'd650066}}},
    '{'{'{25'd150302, -25'd2204423, -25'd551106, -25'd4208444, -25'd300603, -25'd3406835, 25'd400804, 25'd150302, 25'd0}, '{25'd1853719, 25'd3406835, 25'd3356735, 25'd1302614, -25'd751508, 25'd200402, 25'd3807640, 25'd4308645, 25'd601206}, '{25'd2705428, 25'd1503016, -25'd4659348, -25'd2254523, -25'd1102211, 25'd651307, 25'd4509047, -25'd2605227, 25'd3306634}, '{-25'd701407, 25'd501005, 25'd0, -25'd1503016, 25'd551106, 25'd1553116, -25'd3557137, 25'd450905, 25'd4759550}, '{-25'd951910, -25'd400804, -25'd2905830, -25'd4208444, -25'd1202413, 25'd851709, -25'd1503016, -25'd2905830, 25'd250503}, '{25'd2855730, -25'd1553116, -25'd3957941, 25'd601206, 25'd1753518, -25'd1703418, -25'd4108243, 25'd2555127, 25'd4559147}, '{25'd3006031, 25'd1553116, 25'd1703418, -25'd2805629, -25'd4509047, -25'd3106232, -25'd2204423, 25'd1903820, 25'd2204423}, '{25'd2254523, -25'd50101, 25'd1603217, -25'd1452915, 25'd551106, 25'd3657338, -25'd3156333, 25'd1853719, 25'd1903820}, '{-25'd1553116, 25'd601206, 25'd4859751, 25'd4108243, -25'd701407, -25'd901809, -25'd2154322, -25'd100201, 25'd450905}}, '{'{-25'd3507036, 25'd2104222, -25'd501005, 25'd3356735, -25'd350704, 25'd4759550, 25'd1953920, 25'd2054121, 25'd2204423}, '{-25'd200402, -25'd4458946, -25'd1402815, 25'd3156333, 25'd3657338, 25'd5360756, -25'd50101, 25'd1903820, 25'd601206}, '{25'd2004021, -25'd3707439, 25'd701407, -25'd3356735, -25'd3456936, 25'd3957941, 25'd4559147, 25'd1352714, -25'd2154322}, '{25'd100201, 25'd4008042, -25'd5160354, -25'd1953920, -25'd501005, 25'd951910, -25'd2555127, 25'd501005, 25'd4258544}, '{-25'd751508, -25'd3056132, -25'd5060153, -25'd2705428, -25'd5511057, -25'd150302, -25'd751508, 25'd3757539, -25'd3907841}, '{-25'd2204423, -25'd450905, 25'd2204423, 25'd1002010, -25'd6412867, -25'd2755529, -25'd1202413, 25'd2304624, -25'd3657338}, '{25'd3607238, 25'd601206, 25'd250503, 25'd2204423, -25'd551106, 25'd3106232, -25'd3907841, 25'd3356735, -25'd3907841}, '{25'd551106, -25'd2404825, 25'd951910, 25'd2905830, -25'd3056132, 25'd3557137, -25'd3757539, 25'd3306634, -25'd751508}, '{-25'd300603, -25'd1052111, -25'd2905830, 25'd4659348, 25'd4509047, 25'd3406835, 25'd4959952, -25'd3507036, 25'd4058142}}, '{'{-25'd701407, -25'd1452915, -25'd4008042, -25'd2054121, -25'd2354725, 25'd2755529, 25'd300603, 25'd1152312, 25'd751508}, '{25'd2555127, 25'd200402, -25'd250503, 25'd4659348, 25'd2304624, 25'd2004021, 25'd350704, 25'd1402815, -25'd1803619}, '{-25'd100201, 25'd2404825, -25'd1503016, 25'd4859751, -25'd801608, 25'd3607238, 25'd5460957, 25'd4158343, -25'd2104222}, '{25'd1703418, -25'd651307, 25'd3106232, -25'd3006031, 25'd100201, 25'd2555127, 25'd3356735, 25'd1903820, 25'd1953920}, '{25'd250503, -25'd1402815, 25'd4008042, -25'd1903820, -25'd2855730, -25'd3306634, -25'd4008042, 25'd751508, 25'd751508}, '{25'd2054121, -25'd1703418, 25'd350704, 25'd2655328, -25'd5661359, -25'd5410856, -25'd3857740, 25'd1252513, -25'd2204423}, '{25'd2204423, -25'd150302, 25'd2304624, -25'd1753518, -25'd1603217, -25'd2805629, -25'd5661359, -25'd3106232, 25'd2505026}, '{25'd300603, -25'd1402815, 25'd4358745, 25'd2505026, -25'd3056132, 25'd851709, -25'd450905, 25'd1252513, 25'd0}, '{25'd1302614, -25'd651307, -25'd2655328, 25'd350704, 25'd2605227, 25'd1803619, -25'd2505026, -25'd1352714, 25'd3256534}}},
    '{'{'{25'd710201, 25'd3381910, -25'd980754, 25'd845477, -25'd4092111, 25'd3212814, -25'd1116030, 25'd2840804, -25'd777839}, '{25'd4058292, -25'd1690955, 25'd1860050, 25'd1251307, 25'd2468794, 25'd4159749, -25'd4295025, 25'd3517186, -25'd4328844}, '{25'd574925, -25'd1352764, -25'd3043719, 25'd2299699, 25'd4058292, 25'd4159749, 25'd1961508, 25'd1758593, -25'd1183668}, '{-25'd2265879, 25'd2164422, -25'd1521859, 25'd811658, -25'd3178995, 25'd3077538, 25'd3280452, 25'd1589498, 25'd2096784}, '{25'd2773166, 25'd1724774, -25'd2468794, -25'd1116030, -25'd1420402, 25'd3280452, -25'd2773166, 25'd2536432, 25'd1183668}, '{25'd3280452, 25'd3584824, -25'd2942261, -25'd2773166, 25'd2976080, -25'd1420402, 25'd2367337, -25'd2265879, 25'd3821558}, '{-25'd1758593, 25'd2096784, 25'd236734, -25'd2604070, 25'd1758593, -25'd1927688, 25'd169095, 25'd3145176, -25'd202915}, '{25'd2401156, 25'd338191, 25'd676382, 25'd2705528, -25'd2773166, -25'd3821558, -25'd2367337, -25'd1454221, -25'd1488040}, '{25'd913116, 25'd439648, -25'd2333518, -25'd304372, -25'd2062965, -25'd1386583, 25'd338191, -25'd1149849, 25'd2198241}}, '{'{25'd1826231, -25'd2198241, 25'd1454221, -25'd4092111, 25'd642563, 25'd2502613, -25'd135276, 25'd1285126, -25'd439648}, '{25'd0, -25'd2434975, 25'd2908442, 25'd2468794, 25'd0, -25'd744020, 25'd1521859, -25'd2705528, 25'd135276}, '{25'd33819, -25'd574925, -25'd304372, -25'd3686281, -25'd2198241, -25'd3990653, 25'd2062965, -25'd913116, 25'd1082211}, '{-25'd3551005, -25'd1995327, -25'd3551005, 25'd338191, 25'd2570251, -25'd3618643, 25'd1589498, 25'd1217487, -25'd270553}, '{25'd4261206, -25'd1893869, 25'd3246633, 25'd3990653, -25'd101457, -25'd1082211, 25'd2130603, 25'd1082211, -25'd2637889}, '{-25'd2367337, -25'd3111357, 25'd2164422, 25'd3212814, 25'd2468794, -25'd744020, -25'd676382, -25'd1149849, 25'd4227387}, '{-25'd3821558, -25'd1792412, 25'd2367337, 25'd1690955, -25'd1961508, -25'd2029146, -25'd2739347, -25'd1454221, -25'd3517186}, '{-25'd3652462, -25'd2299699, -25'd236734, 25'd2637889, -25'd3348091, 25'd2130603, 25'd1318945, -25'd2806985, -25'd2908442}, '{-25'd2401156, -25'd744020, 25'd608744, -25'd3483367, -25'd3753920, -25'd2265879, -25'd1318945, -25'd2130603, 25'd2570251}}, '{'{25'd3212814, 25'd3483367, -25'd1961508, 25'd1657136, 25'd2434975, 25'd2806985, 25'd1116030, 25'd2570251, -25'd676382}, '{-25'd642563, 25'd2671709, -25'd1555678, 25'd33819, -25'd2198241, 25'd202915, -25'd2029146, 25'd3923015, -25'd3145176}, '{-25'd3178995, -25'd1217487, 25'd3990653, -25'd3314271, -25'd811658, -25'd2130603, -25'd2198241, -25'd1555678, 25'd3314271}, '{-25'd338191, 25'd1251307, -25'd3720101, -25'd2096784, 25'd744020, 25'd3618643, -25'd980754, 25'd1285126, 25'd2029146}, '{-25'd1420402, -25'd1318945, -25'd135276, 25'd2773166, -25'd2401156, -25'd1488040, 25'd2671709, -25'd777839, 25'd1995327}, '{-25'd372010, -25'd2536432, -25'd2671709, -25'd2705528, 25'd1217487, -25'd1251307, 25'd4227387, 25'd3889196, 25'd4024472}, '{-25'd3889196, 25'd2265879, 25'd2401156, 25'd2029146, -25'd4058292, 25'd3449548, 25'd4024472, -25'd3956834, -25'd541106}, '{25'd270553, -25'd3212814, 25'd2739347, -25'd67638, 25'd3348091, 25'd2908442, -25'd1860050, -25'd3889196, 25'd439648}, '{25'd1792412, 25'd3009900, 25'd3111357, -25'd1589498, 25'd1724774, 25'd1758593, 25'd3821558, 25'd2130603, -25'd338191}}},
    '{'{'{-25'd2759998, -25'd1433765, -25'd394285, -25'd3512725, 25'd2903374, -25'd3763634, -25'd4444672, -25'd501818, 25'd2150648}, '{-25'd3225972, -25'd215065, -25'd2150648, -25'd465974, 25'd3942854, 25'd609350, -25'd3584413, -25'd2294024, -25'd2294024}, '{-25'd1612986, 25'd896103, 25'd609350, 25'd3799478, 25'd3512725, 25'd3727789, -25'd4193763, -25'd681038, 25'd1863895}, '{-25'd2903374, -25'd2688310, 25'd3261816, 25'd2401557, 25'd1147012, 25'd358441, 25'd3154283, -25'd286753, 25'd716883}, '{25'd3978698, 25'd143377, 25'd4157919, 25'd3835322, 25'd465974, 25'd3441036, 25'd215065, 25'd824415, -25'd4193763}, '{-25'd3835322, 25'd967791, -25'd967791, 25'd1147012, -25'd2867530, -25'd1469609, -25'd501818, 25'd4050387, -25'd1720518}, '{-25'd2759998, 25'd1218700, 25'd1362077, 25'd3297660, 25'd3476881, 25'd3548569, -25'd2329868, -25'd3441036, -25'd3297660}, '{25'd2222336, -25'd1505453, 25'd1577142, -25'd1469609, 25'd2580777, -25'd1899739, 25'd3548569, 25'd1720518, 25'd3046751}, '{-25'd3656101, 25'd2688310, 25'd4229607, 25'd1075324, -25'd2222336, -25'd3799478, -25'd3190127, -25'd2258180, 25'd2150648}}, '{'{25'd1397921, 25'd1326233, 25'd1218700, 25'd215065, 25'd1505453, -25'd3261816, 25'd1541298, -25'd931947, -25'd3441036}, '{-25'd250909, 25'd394285, 25'd215065, 25'd3727789, 25'd250909, 25'd3046751, 25'd1720518, -25'd3333504, 25'd3691945}, '{-25'd286753, -25'd1075324, 25'd1720518, 25'd1147012, -25'd2759998, 25'd716883, 25'd2329868, -25'd2509089, -25'd2258180}, '{25'd3942854, -25'd3691945, 25'd573506, -25'd3046751, 25'd2509089, -25'd2222336, 25'd2867530, -25'd4050387, -25'd2473245}, '{25'd3978698, -25'd4444672, 25'd2616621, -25'd2867530, -25'd1505453, -25'd1541298, -25'd2186492, 25'd1720518, -25'd967791}, '{25'd2616621, -25'd3190127, 25'd1182856, 25'd3548569, -25'd2652466, -25'd967791, 25'd967791, 25'd3190127, 25'd1182856}, '{-25'd143377, -25'd2078959, 25'd3656101, -25'd1577142, -25'd179221, -25'd3010907, -25'd1541298, 25'd2078959, -25'd71688}, '{25'd3154283, 25'd3907010, -25'd824415, 25'd2939219, -25'd752727, -25'd2616621, -25'd4552204, -25'd2043115, -25'd3476881}, '{-25'd3620257, -25'd3691945, -25'd501818, 25'd931947, -25'd1182856, 25'd286753, 25'd3548569, -25'd3190127, 25'd2365713}}, '{'{25'd2258180, -25'd860259, 25'd1935583, 25'd1290389, 25'd2867530, -25'd4086231, -25'd1863895, -25'd573506, 25'd2867530}, '{-25'd3871166, 25'd1577142, 25'd2150648, 25'd3584413, -25'd4408828, 25'd430130, -25'd394285, 25'd3871166, -25'd2365713}, '{25'd179221, 25'd322597, -25'd3297660, -25'd1505453, 25'd1433765, 25'd2329868, 25'd2258180, -25'd3046751, 25'd860259}, '{-25'd2437401, -25'd3154283, 25'd1147012, -25'd3978698, 25'd215065, -25'd430130, -25'd4086231, -25'd4265451, 25'd1147012}, '{25'd3010907, -25'd1541298, 25'd2544933, 25'd1039480, -25'd1684674, 25'd465974, 25'd3799478, 25'd1612986, -25'd4337140}, '{-25'd4122075, 25'd2186492, -25'd2329868, 25'd2580777, 25'd3656101, -25'd967791, 25'd967791, 25'd1290389, 25'd3691945}, '{-25'd3297660, -25'd4157919, -25'd430130, 25'd3441036, -25'd2867530, 25'd107532, 25'd2724154, 25'd2258180, 25'd4014542}, '{25'd1075324, 25'd3154283, 25'd537662, -25'd3046751, -25'd931947, -25'd1863895, 25'd1648830, 25'd3548569, 25'd35844}, '{-25'd3154283, -25'd1577142, 25'd2007271, -25'd1433765, -25'd4122075, -25'd3010907, 25'd2007271, 25'd3691945, 25'd3942854}}},
    '{'{'{25'd4172062, 25'd1772203, 25'd443051, 25'd3544406, -25'd3729011, 25'd1218390, 25'd2695226, 25'd3950536, 25'd2953672}, '{-25'd1587599, 25'd516893, -25'd3544406, 25'd332288, -25'd1919887, -25'd36921, -25'd2879830, 25'd258446, -25'd2879830}, '{-25'd2916751, -25'd1624520, 25'd2436779, 25'd3692090, -25'd443051, 25'd1181469, -25'd1661441, 25'd886102, 25'd295367}, '{25'd1181469, 25'd4393587, 25'd775339, 25'd2067570, 25'd3913615, -25'd36921, 25'd701497, 25'd2916751, -25'd3064435}, '{-25'd3802853, 25'd443051, -25'd1439915, 25'd2178333, -25'd3729011, 25'd4504350, 25'd110763, -25'd553814, -25'd923023}, '{25'd2695226, 25'd4135141, 25'd221525, -25'd1550678, -25'd2916751, 25'd4615113, 25'd553814, 25'd2510621, 25'd3322881}, '{-25'd2547542, -25'd3359802, 25'd2879830, 25'd2326017, -25'd479972, 25'd1772203, -25'd2289096, 25'd3396723, -25'd2030650}, '{25'd2916751, -25'd1144548, 25'd2326017, -25'd959943, -25'd36921, 25'd2879830, -25'd3285960, -25'd2547542, -25'd2621384}, '{25'd1698361, -25'd3913615, 25'd2990593, -25'd3950536, -25'd2990593, -25'd3322881, 25'd2547542, 25'd3802853, 25'd4024378}}, '{'{25'd4098220, 25'd4393587, -25'd258446, 25'd1476836, 25'd1292232, 25'd3359802, 25'd1218390, -25'd2584463, 25'd3802853}, '{-25'd73842, -25'd553814, 25'd4061299, -25'd3396723, -25'd3876695, -25'd3433644, -25'd2289096, -25'd1366073, -25'd2916751}, '{-25'd1070706, 25'd2842909, 25'd3692090, 25'd4245904, -25'd3138277, 25'd3249039, -25'd3692090, -25'd3507486, -25'd1882966}, '{25'd2695226, 25'd886102, -25'd2621384, 25'd2141412, -25'd443051, -25'd2215254, -25'd1882966, -25'd1919887, 25'd2473700}, '{25'd1070706, -25'd1550678, -25'd2362938, -25'd2473700, -25'd2141412, 25'd4541271, 25'd3249039, 25'd3027514, -25'd110763}, '{25'd2399859, -25'd1329152, -25'd738418, -25'd1513757, 25'd1476836, -25'd2326017, 25'd4282824, 25'd73842, -25'd886102}, '{25'd1587599, 25'd3027514, -25'd1366073, -25'd3655169, 25'd1218390, 25'd258446, -25'd2436779, 25'd295367, -25'd1439915}, '{25'd443051, 25'd332288, -25'd443051, 25'd2067570, 25'd4135141, -25'd3285960, -25'd2658305, 25'd3913615, 25'd2547542}, '{-25'd2362938, -25'd406130, 25'd3729011, -25'd4024378, 25'd2067570, 25'd3507486, -25'd3765932, -25'd1476836, -25'd3470565}}, '{'{-25'd738418, 25'd2879830, 25'd3212118, -25'd1846045, -25'd3729011, 25'd4393587, -25'd775339, 25'd1846045, -25'd3433644}, '{25'd3433644, 25'd923023, 25'd1809124, 25'd258446, -25'd959943, 25'd1956808, 25'd4393587, 25'd4135141, 25'd2547542}, '{25'd775339, -25'd3396723, -25'd2732147, -25'd3285960, 25'd4393587, -25'd443051, 25'd1366073, 25'd479972, 25'd701497}, '{-25'd1735282, 25'd4430508, 25'd1550678, 25'd3876695, 25'd2030650, 25'd2805988, -25'd2326017, 25'd3064435, -25'd1513757}, '{25'd4541271, -25'd1033785, 25'd1402994, -25'd1144548, -25'd1218390, -25'd3618248, -25'd3802853, 25'd3101356, -25'd1070706}, '{-25'd2547542, 25'd886102, 25'd406130, 25'd4688954, 25'd147684, 25'd2326017, -25'd1144548, 25'd2030650, 25'd775339}, '{-25'd2289096, 25'd258446, -25'd812260, 25'd738418, 25'd4504350, 25'd2805988, -25'd701497, -25'd2141412, -25'd1698361}, '{-25'd627655, 25'd2030650, 25'd3729011, -25'd1476836, 25'd4430508, 25'd36921, 25'd2067570, -25'd2067570, 25'd4319745}, '{-25'd2399859, -25'd221525, 25'd443051, 25'd258446, -25'd1772203, -25'd3618248, 25'd1772203, -25'd2067570, 25'd3987457}}},
    '{'{'{-25'd2922014, -25'd3146785, 25'd2060395, -25'd2847091, -25'd1123852, 25'd2397550, 25'd1498469, 25'd1461007, -25'd1236237}, '{-25'd711773, 25'd74923, 25'd1535931, 25'd1535931, 25'd3746172, 25'd2322627, -25'd3146785, 25'd0, -25'd1798163}, '{25'd749234, -25'd3821096, 25'd1948010, 25'd1236237, 25'd2884553, 25'd3896019, -25'd2210242, -25'd4045866, 25'd2884553}, '{25'd1873086, 25'd3521402, 25'd1573392, 25'd1386084, 25'd974005, -25'd599388, 25'd1835624, -25'd3409017, 25'd561926}, '{25'd4308098, -25'd187309, 25'd749234, 25'd3259170, 25'd3221708, 25'd3184246, -25'd2285165, 25'd899081, -25'd2996938}, '{-25'd3371555, 25'd3708711, 25'd2397550, -25'd3783634, 25'd899081, -25'd449541, -25'd4795100, -25'd1273699, -25'd2659782}, '{25'd974005, -25'd2734706, -25'd1311160, 25'd1011467, -25'd37462, -25'd1461007, 25'd2397550, -25'd3858557, 25'd2210242}, '{-25'd3296632, -25'd936543, 25'd1685778, 25'd1573392, 25'd2697244, -25'd4345560, 25'd1348622, 25'd1685778, -25'd2060395}, '{-25'd2884553, -25'd4158251, -25'd3071861, 25'd3858557, -25'd4195713, -25'd3296632, -25'd3970943, -25'd1535931, 25'd2022933}}, '{'{25'd2809629, -25'd487002, 25'd4158251, 25'd936543, 25'd1723239, -25'd1535931, 25'd3858557, 25'd187309, 25'd2210242}, '{-25'd3783634, -25'd2809629, 25'd4158251, 25'd3970943, -25'd824158, 25'd2097856, -25'd1685778, -25'd3896019, 25'd786696}, '{-25'd2547397, 25'd1123852, 25'd1985471, -25'd3371555, 25'd3633787, -25'd2547397, 25'd3296632, -25'd2210242, 25'd1236237}, '{25'd1386084, -25'd1498469, 25'd2097856, 25'd4158251, 25'd2622321, 25'd2060395, 25'd3184246, -25'd1648316, -25'd1048928}, '{25'd936543, -25'd3409017, 25'd1198775, -25'd3708711, 25'd1161313, -25'd3970943, -25'd2772167, 25'd2734706, -25'd1011467}, '{25'd3596325, -25'd2547397, -25'd4495407, -25'd449541, -25'd449541, 25'd412079, -25'd4195713, 25'd3446478, -25'd2809629}, '{25'd74923, -25'd2172780, -25'd1011467, -25'd1048928, 25'd299694, 25'd636849, 25'd936543, -25'd749234, -25'd2772167}, '{25'd3109323, 25'd3933481, 25'd487002, 25'd974005, -25'd3071861, 25'd599388, -25'd1348622, -25'd3034400, 25'd1498469}, '{-25'd3596325, 25'd2135318, -25'd2772167, 25'd1348622, -25'd1123852, 25'd1798163, -25'd224770, -25'd2509935, -25'd3071861}}, '{'{-25'd1161313, 25'd936543, -25'd2322627, -25'd3146785, 25'd3221708, -25'd3783634, -25'd1535931, 25'd3146785, -25'd2360089}, '{25'd3708711, 25'd3521402, -25'd599388, 25'd3146785, -25'd3970943, -25'd2996938, -25'd3071861, -25'd1423545, 25'd149847}, '{25'd2172780, 25'd2584859, -25'd4645254, -25'd4645254, 25'd1161313, 25'd1423545, -25'd187309, -25'd3596325, 25'd3409017}, '{25'd449541, -25'd3671249, -25'd636849, 25'd1760701, 25'd1535931, -25'd4083328, -25'd2697244, 25'd1985471, -25'd4195713}, '{25'd936543, 25'd2247703, 25'd3371555, 25'd561926, -25'd37462, 25'd299694, -25'd4270636, -25'd3184246, 25'd3334093}, '{-25'd2509935, 25'd1910548, 25'd3109323, -25'd2472474, 25'd0, -25'd4757639, -25'd1423545, 25'd2472474, 25'd711773}, '{-25'd4420483, 25'd3259170, -25'd749234, -25'd4158251, -25'd74923, 25'd3221708, -25'd4795100, 25'd1461007, 25'd861620}, '{-25'd2547397, 25'd1311160, -25'd3334093, 25'd74923, -25'd3446478, 25'd1461007, 25'd2772167, -25'd4795100, -25'd4795100}, '{25'd2622321, -25'd2547397, -25'd3896019, 25'd2959476, -25'd4795100, 25'd1648316, 25'd711773, -25'd3558864, -25'd2097856}}},
    '{'{'{25'd3580109, -25'd1716991, -25'd2739879, -25'd73063, 25'd730634, 25'd3762768, 25'd730634, 25'd1315142, 25'd3945426}, '{25'd4274212, -25'd3324387, 25'd3397450, 25'd4128085, -25'd2995601, -25'd949825, -25'd694103, -25'd4091553, -25'd219190}, '{25'd1607396, -25'd3689704, 25'd2155372, -25'd1899650, 25'd4164617, 25'd2338030, 25'd73063, 25'd0, -25'd3762768}, '{-25'd3616641, 25'd1570864, 25'd2009245, -25'd2995601, 25'd2009245, 25'd1607396, 25'd2995601, 25'd401849, 25'd1169015}, '{25'd949825, -25'd2703348, -25'd255722, 25'd4493402, -25'd3433982, 25'd2520689, 25'd2264967, 25'd4128085, 25'd986357}, '{-25'd3981958, -25'd4237680, 25'd255722, -25'd2959070, 25'd986357, 25'd1424737, -25'd986357, 25'd2593752, 25'd1790054}, '{-25'd146127, -25'd2703348, -25'd3872363, -25'd1753523, 25'd986357, -25'd2338030, -25'd3105197, 25'd3214792, 25'd4128085}, '{25'd4420339, 25'd3141728, 25'd365317, 25'd840230, -25'd3251323, -25'd3141728, -25'd3178260, 25'd3068665, -25'd3689704}, '{-25'd1278610, -25'd1972713, -25'd2776411, -25'd2045777, -25'd2520689, -25'd2484157, 25'd1534332, 25'd876761, -25'd3580109}}, '{'{-25'd2849474, -25'd2082308, 25'd2593752, -25'd2812943, -25'd2995601, 25'd2155372, 25'd3908894, 25'd621039, -25'd2082308}, '{-25'd3324387, -25'd292254, -25'd3726236, -25'd3214792, -25'd2886006, 25'd4529934, -25'd182659, 25'd3799299, 25'd4018490}, '{25'd2922538, -25'd3507046, 25'd1716991, -25'd2264967, 25'd2228435, -25'd3543577, -25'd3507046, -25'd3141728, -25'd1534332}, '{-25'd182659, 25'd3981958, 25'd949825, 25'd621039, -25'd2776411, -25'd1497801, 25'd2959070, -25'd1570864, -25'd3762768}, '{25'd3872363, -25'd2338030, -25'd4420339, 25'd255722, 25'd1132483, 25'd511444, 25'd1022888, -25'd2995601, -25'd3945426}, '{25'd1022888, -25'd2959070, 25'd2009245, -25'd2557221, -25'd4456870, 25'd1461269, 25'd730634, -25'd2374562, -25'd2630284}, '{-25'd1716991, 25'd1972713, -25'd182659, -25'd2338030, -25'd4493402, 25'd2191903, -25'd3908894, 25'd3835831, -25'd146127}, '{25'd1899650, -25'd182659, 25'd3616641, -25'd986357, -25'd1059420, 25'd767166, 25'd4639529, -25'd3507046, -25'd584508}, '{25'd2264967, 25'd3835831, -25'd3507046, 25'd4566466, 25'd3908894, 25'd4164617, 25'd1863118, 25'd4639529, 25'd4566466}}, '{'{25'd2118840, -25'd3835831, -25'd2118840, -25'd2922538, 25'd4237680, -25'd3653172, 25'd1716991, -25'd1205547, -25'd1716991}, '{-25'd1826586, 25'd4383807, -25'd3032133, 25'd146127, 25'd2301499, 25'd2520689, -25'd3178260, 25'd3872363, 25'd584508}, '{25'd2264967, 25'd2301499, -25'd1570864, -25'd474912, 25'd438381, 25'd474912, -25'd3068665, -25'd3653172, 25'd2520689}, '{25'd3287855, 25'd1059420, -25'd986357, -25'd4310743, -25'd2922538, 25'd474912, -25'd1936181, 25'd3178260, 25'd2155372}, '{25'd2045777, -25'd438381, 25'd3799299, 25'd2593752, -25'd1936181, 25'd1570864, 25'd474912, 25'd2082308, -25'd3397450}, '{-25'd1351674, 25'd3908894, 25'd36532, -25'd1388206, -25'd3141728, -25'd3178260, -25'd2630284, -25'd4201148, 25'd4274212}, '{-25'd3507046, 25'd255722, -25'd3068665, 25'd3835831, -25'd3068665, 25'd2922538, 25'd1534332, -25'd146127, 25'd803698}, '{25'd3908894, -25'd621039, 25'd1132483, -25'd1022888, -25'd1972713, -25'd2849474, -25'd1936181, 25'd3835831, 25'd3251323}, '{-25'd2703348, -25'd2082308, 25'd2082308, 25'd438381, -25'd2374562, -25'd1351674, 25'd1716991, 25'd4639529, 25'd1497801}}},
    '{'{'{25'd2967700, -25'd1951365, -25'd894375, -25'd3496195, 25'd3089661, -25'd487841, -25'd3130314, 25'd3130314, 25'd4187303}, '{-25'd2235939, 25'd1748097, -25'd3211621, 25'd4309264, 25'd2967700, 25'd2520513, -25'd3618155, -25'd894375, 25'd447188}, '{25'd243921, -25'd2439206, 25'd2805087, -25'd1707444, -25'd447188, 25'd1138296, -25'd2317245, -25'd569148, -25'd975682}, '{25'd2357899, 25'd3577502, -25'd2683126, -25'd528495, 25'd1016336, 25'd650455, -25'd121960, -25'd2845740, 25'd40653}, '{25'd1463523, 25'd3049007, -25'd3130314, -25'd1138296, 25'd1219603, 25'd1138296, 25'd731762, -25'd650455, 25'd1951365}, '{-25'd1138296, 25'd3902729, 25'd3577502, 25'd4756451, 25'd650455, -25'd162614, -25'd1829404, -25'd2886393, -25'd3536848}, '{25'd528495, 25'd935029, -25'd3089661, 25'd4471877, 25'd1260256, 25'd1260256, 25'd3292928, -25'd1341563, -25'd40653}, '{-25'd3292928, 25'd3984036, 25'd2398552, 25'd4105996, -25'd894375, 25'd4065343, -25'd406534, 25'd2154632, 25'd406534}, '{25'd1951365, -25'd1788751, -25'd2479859, 25'd1219603, 25'd203267, 25'd2886393, 25'd2886393, 25'd2317245, -25'd1788751}}, '{'{-25'd3577502, -25'd691108, -25'd935029, -25'd2886393, -25'd1829404, 25'd4309264, -25'd40653, 25'd1260256, 25'd3292928}, '{-25'd3089661, 25'd2195285, -25'd1422870, 25'd772415, -25'd1016336, 25'd1870058, -25'd1666791, -25'd2805087, -25'd3292928}, '{25'd121960, 25'd731762, -25'd2479859, 25'd3902729, 25'd691108, -25'd3374235, 25'd487841, 25'd1585484, -25'd1300910}, '{25'd1544830, 25'd650455, -25'd3699462, 25'd4553184, 25'd284574, -25'd2886393, -25'd2317245, 25'd4227957, 25'd1382217}, '{25'd3618155, 25'd2927047, 25'd1382217, 25'd609801, 25'd1748097, -25'd935029, -25'd1626137, 25'd4431224, -25'd731762}, '{25'd3943383, 25'd81307, 25'd813069, 25'd203267, -25'd1260256, -25'd81307, 25'd2561166, 25'd3699462, 25'd1016336}, '{-25'd2479859, -25'd731762, -25'd1138296, 25'd1748097, 25'd121960, -25'd2683126, -25'd2927047, 25'd2439206, 25'd2561166}, '{25'd3414888, 25'd2073325, 25'd691108, 25'd5081679, 25'd5162986, 25'd3618155, 25'd3496195, 25'd3943383, -25'd1992018}, '{-25'd1951365, 25'd3374235, 25'd2479859, 25'd3333581, 25'd569148, 25'd1829404, 25'd365881, 25'd1504177, 25'd853722}}, '{'{25'd3049007, -25'd3089661, 25'd3049007, -25'd1626137, 25'd243921, -25'd3618155, 25'd1910711, 25'd2845740, -25'd3943383}, '{-25'd3618155, -25'd813069, 25'd365881, -25'd2479859, -25'd3455542, -25'd3658809, -25'd4024690, 25'd1829404, -25'd2601819}, '{-25'd1463523, 25'd447188, 25'd2967700, -25'd3902729, 25'd243921, -25'd2764433, -25'd1504177, -25'd813069, 25'd447188}, '{25'd1666791, -25'd2073325, -25'd4593838, 25'd2439206, 25'd3658809, -25'd2317245, 25'd162614, 25'd731762, 25'd365881}, '{-25'd3130314, -25'd284574, 25'd1829404, -25'd3699462, 25'd4349917, 25'd1382217, -25'd81307, -25'd487841, 25'd691108}, '{-25'd528495, 25'd162614, -25'd3862076, -25'd3862076, 25'd2317245, 25'd4593838, 25'd528495, -25'd81307, -25'd243921}, '{25'd2927047, -25'd1585484, 25'd3455542, -25'd3577502, 25'd2561166, -25'd731762, 25'd3740116, -25'd4187303, -25'd3902729}, '{-25'd365881, 25'd406534, 25'd4187303, 25'd691108, 25'd1788751, -25'd3496195, 25'd894375, 25'd1666791, 25'd81307}, '{-25'd243921, -25'd3618155, -25'd1504177, -25'd3984036, 25'd1504177, 25'd3862076, 25'd3211621, -25'd1748097, -25'd2642473}}},
    '{'{'{-25'd3460638, -25'd3142824, 25'd1412505, -25'd3813764, -25'd953441, 25'd353126, -25'd2577822, 25'd211876, 25'd882816}, '{-25'd3672513, -25'd3743139, 25'd4272828, -25'd176563, -25'd247188, -25'd3178136, -25'd1271255, -25'd2683760, 25'd1765631}, '{25'd2825010, -25'd600315, 25'd1483130, -25'd776878, -25'd1024066, -25'd1412505, 25'd3390012, -25'd70625, 25'd2930948}, '{-25'd600315, -25'd388439, -25'd1765631, 25'd317814, 25'd1271255, 25'd2648447, 25'd1800944, 25'd3178136, 25'd2083445}, '{-25'd741565, 25'd4378766, -25'd1942195, 25'd105938, -25'd3990327, 25'd1200629, -25'd3425325, 25'd635627, -25'd1341880}, '{25'd2012820, 25'd847503, -25'd1624381, -25'd2330633, -25'd2754385, 25'd2189383, 25'd1836257, -25'd3248762, -25'd459064}, '{-25'd918128, -25'd3425325, 25'd706253, 25'd4484704, 25'd282501, 25'd2118758, -25'd3778451, 25'd1130004, 25'd3566575}, '{25'd3319387, -25'd635627, 25'd3107511, 25'd2754385, 25'd3142824, -25'd247188, 25'd3707826, -25'd3107511, 25'd2118758}, '{25'd1765631, 25'd3142824, 25'd3142824, -25'd2260008, -25'd918128, -25'd2401259, 25'd4414078, 25'd4378766, 25'd1518443}}, '{'{-25'd1624381, 25'd3390012, -25'd2154070, 25'd2471884, -25'd1377192, -25'd1412505, -25'd423752, 25'd3213449, 25'd3495950}, '{-25'd953441, 25'd282501, 25'd600315, -25'd2224696, -25'd2507197, 25'd353126, -25'd741565, -25'd4060952, -25'd1094691}, '{-25'd1836257, 25'd282501, 25'd247188, -25'd2295321, 25'd3036886, -25'd2648447, -25'd3036886, -25'd3955014, 25'd3319387}, '{25'd2401259, 25'd1659694, 25'd4484704, 25'd3001573, -25'd2189383, -25'd1589068, -25'd3990327, 25'd2507197, 25'd2154070}, '{-25'd2154070, 25'd3955014, -25'd1377192, 25'd459064, 25'd4060952, -25'd3248762, 25'd3390012, 25'd70625, -25'd918128}, '{-25'd2118758, 25'd459064, 25'd3919702, -25'd3425325, 25'd1200629, 25'd1730319, -25'd3001573, 25'd1589068, -25'd3990327}, '{25'd2719072, 25'd741565, -25'd2365946, -25'd2224696, 25'd176563, -25'd3001573, -25'd2189383, -25'd2224696, -25'd70625}, '{-25'd3707826, 25'd2719072, 25'd1765631, -25'd2860323, -25'd2789698, -25'd4166890, 25'd35313, -25'd2330633, 25'd247188}, '{-25'd2083445, 25'd2754385, -25'd2436571, 25'd353126, 25'd3955014, 25'd2436571, 25'd2789698, 25'd882816, -25'd706253}}, '{'{25'd2401259, 25'd2966261, 25'd317814, -25'd3390012, 25'd2471884, 25'd1483130, 25'd1024066, -25'd353126, 25'd1977507}, '{-25'd2189383, -25'd2012820, 25'd353126, -25'd247188, -25'd1659694, 25'd3178136, 25'd1094691, 25'd2224696, -25'd2012820}, '{-25'd1165317, -25'd3248762, -25'd2895635, -25'd4025640, 25'd4484704, -25'd1659694, -25'd2825010, 25'd2542509, 25'd211876}, '{-25'd3284074, 25'd600315, 25'd3990327, 25'd3178136, 25'd2542509, 25'd2895635, -25'd1094691, -25'd3566575, -25'd2507197}, '{-25'd529689, -25'd3213449, 25'd1730319, -25'd1695006, -25'd3001573, 25'd4414078, 25'd2436571, 25'd2648447, -25'd3566575}, '{25'd2189383, -25'd2260008, 25'd176563, 25'd1200629, -25'd2295321, -25'd2825010, 25'd670940, -25'd3778451, -25'd4237515}, '{-25'd1200629, -25'd2224696, 25'd953441, 25'd3495950, -25'd2471884, 25'd2613134, 25'd882816, 25'd3849076, -25'd1906882}, '{25'd3707826, -25'd423752, 25'd882816, -25'd918128, 25'd3813764, 25'd3390012, 25'd882816, 25'd211876, -25'd4237515}, '{25'd2295321, -25'd4202203, -25'd353126, -25'd2966261, 25'd2189383, 25'd3284074, -25'd282501, -25'd1059379, 25'd3284074}}},
    '{'{'{25'd2216798, 25'd1125993, -25'd2639045, 25'd4152097, 25'd1935300, 25'd2287172, -25'd2639045, 25'd3166854, 25'd4328034}, '{25'd1618614, -25'd1090805, -25'd1794551, 25'd2533483, -25'd3518727, -25'd1090805, -25'd1055618, 25'd2885356, 25'd2498296}, '{25'd4292846, -25'd2850169, -25'd2603858, 25'd3237228, 25'd1548240, -25'd1794551, 25'd4011348, 25'd1196367, -25'd1090805}, '{25'd809307, -25'd562996, 25'd2568670, 25'd1020431, -25'd2392734, -25'd3659476, 25'd1794551, -25'd1688989, -25'd4257659}, '{25'd2040861, 25'd3096479, -25'd562996, 25'd1337116, -25'd3448352, -25'd2076049, 25'd1583427, 25'd1090805, 25'd3940974}, '{-25'd70375, -25'd3659476, -25'd211124, 25'd105562, 25'd3131667, 25'd844494, -25'd598184, 25'd4116910, -25'd281498}, '{-25'd457434, -25'd3976161, 25'd4433596, -25'd2040861, 25'd3624288, 25'd2955730, -25'd3342790, -25'd1653801, -25'd1161180}, '{25'd1337116, -25'd1125993, 25'd3377978, -25'd703745, -25'd3518727, 25'd1442678, -25'd2885356, -25'd1688989, -25'd2568670}, '{-25'd844494, 25'd3518727, 25'd1829738, -25'd351873, -25'd2040861, -25'd2322360, 25'd3448352, -25'd3553914, 25'd1442678}}, '{'{-25'd3377978, 25'd70375, 25'd316685, -25'd809307, 25'd1477865, -25'd1583427, 25'd2814981, 25'd3342790, -25'd2498296}, '{25'd2463109, 25'd1935300, -25'd2885356, 25'd527809, 25'd4328034, 25'd2392734, 25'd2463109, 25'd4081723, 25'd457434}, '{25'd1688989, 25'd1724176, -25'd3659476, 25'd2533483, -25'd1301929, -25'd1864925, 25'd2639045, 25'd3518727, 25'd1759363}, '{25'd1759363, -25'd3377978, 25'd3659476, -25'd2779794, -25'd1618614, 25'd4468783, 25'd1055618, 25'd4433596, -25'd2181610}, '{-25'd211124, 25'd35187, 25'd4187285, 25'd2357547, -25'd1618614, 25'd3729850, -25'd3589101, -25'd1090805, -25'd492622}, '{-25'd3377978, -25'd70375, 25'd4152097, -25'd1970487, -25'd3272416, 25'd668558, 25'd1196367, -25'd2076049, -25'd422247}, '{25'd2639045, 25'd3166854, -25'd351873, 25'd1583427, 25'd3518727, -25'd387060, -25'd35187, -25'd4152097, -25'd2427921}, '{25'd3272416, -25'd1196367, 25'd2674232, -25'd140749, 25'd3202041, -25'd2005674, 25'd985243, 25'd2322360, -25'd1618614}, '{-25'd2251985, 25'd492622, 25'd1407491, -25'd2111236, -25'd2850169, -25'd4116910, 25'd140749, 25'd774120, 25'd2392734}}, '{'{25'd1513052, -25'd3659476, 25'd2146423, -25'd1829738, 25'd3413165, 25'd1301929, 25'd4011348, 25'd1301929, -25'd3272416}, '{-25'd3342790, 25'd4222472, 25'd175936, 25'd1794551, -25'd3342790, -25'd2744607, -25'd1442678, 25'd1759363, -25'd457434}, '{25'd4222472, -25'd1583427, 25'd985243, 25'd3413165, 25'd2850169, 25'd422247, 25'd1688989, 25'd2322360, 25'd3940974}, '{25'd4363221, 25'd1688989, -25'd527809, -25'd950056, 25'd3624288, 25'd1548240, 25'd4257659, -25'd1618614, -25'd2955730}, '{25'd1231554, 25'd1477865, 25'd3096479, 25'd457434, 25'd1829738, -25'd562996, -25'd2568670, -25'd1231554, -25'd703745}, '{-25'd3624288, -25'd3342790, 25'd3131667, 25'd4363221, 25'd387060, -25'd2885356, 25'd4011348, 25'd598184, 25'd4292846}, '{-25'd3800225, 25'd774120, 25'd1055618, 25'd2463109, -25'd1759363, 25'd1724176, 25'd4468783, 25'd1618614, 25'd3131667}, '{25'd1513052, -25'd35187, -25'd2955730, 25'd3377978, -25'd1266742, 25'd3342790, 25'd2990918, 25'd2463109, 25'd2955730}, '{-25'd387060, -25'd4116910, -25'd1864925, -25'd70375, 25'd3659476, -25'd3659476, 25'd3800225, -25'd2357547, 25'd1020431}}},
    '{'{'{25'd1927072, 25'd1745273, -25'd2363391, 25'd763557, 25'd109080, 25'd836277, 25'd2945148, 25'd3054228, 25'd945356}, '{25'd1490754, -25'd3781425, 25'd472678, -25'd4145024, -25'd1854353, 25'd1272595, 25'd1308955, 25'd1636194, 25'd36360}, '{-25'd1636194, 25'd3599626, 25'd72720, 25'd3563266, -25'd581758, -25'd1672553, -25'd2072512, -25'd2108872, 25'd2690629}, '{25'd1272595, -25'd4363183, 25'd36360, 25'd3490546, 25'd3090588, -25'd981716, -25'd3381467, 25'd2036152, 25'd1418034}, '{-25'd727197, 25'd1527114, 25'd2872429, -25'd1745273, -25'd1272595, 25'd2945148, 25'd1199875, -25'd945356, 25'd1454394}, '{-25'd3890505, 25'd2654270, -25'd1454394, 25'd1854353, -25'd145439, -25'd4363183, -25'd2072512, -25'd2108872, -25'd2181591}, '{-25'd872637, 25'd2836069, 25'd1708913, 25'd327239, 25'd1345315, -25'd3890505, -25'd2581550, 25'd1345315, 25'd1018076}, '{-25'd3163308, -25'd690837, -25'd4654062, -25'd1090796, 25'd327239, 25'd4399543, 25'd4326823, 25'd2981508, -25'd2363391}, '{-25'd2508830, -25'd1272595, -25'd4654062, -25'd436318, -25'd1963432, 25'd4108664, 25'd763557, 25'd2763349, 25'd436318}}, '{'{25'd2799709, 25'd2981508, -25'd2436110, 25'd2436110, 25'd3454186, -25'd4435903, 25'd981716, 25'd1490754, 25'd1490754}, '{-25'd836277, -25'd2545190, -25'd2690629, -25'd4108664, -25'd3817785, 25'd4145024, 25'd2472470, -25'd2472470, 25'd509038}, '{-25'd1817993, 25'd3963224, -25'd1963432, -25'd545398, 25'd3054228, -25'd1999792, -25'd727197, -25'd1090796, -25'd1708913}, '{-25'd1672553, -25'd3454186, 25'd363599, -25'd4326823, -25'd3635986, 25'd908996, -25'd1090796, -25'd2726989, -25'd3926865}, '{25'd2399751, -25'd1563474, 25'd1418034, -25'd4654062, -25'd3272387, -25'd908996, 25'd2290671, -25'd2145232, 25'd3599626}, '{25'd2908789, -25'd2217951, -25'd3236027, -25'd2508830, 25'd290879, -25'd1745273, -25'd3963224, 25'd2581550, 25'd3490546}, '{-25'd2763349, -25'd2763349, -25'd4654062, 25'd945356, 25'd3199667, 25'd72720, -25'd2836069, 25'd2290671, 25'd2508830}, '{25'd3272387, -25'd4254103, -25'd218159, -25'd4654062, 25'd1236235, 25'd3126948, 25'd4581342, 25'd3345107, 25'd763557}, '{25'd1817993, 25'd3054228, 25'd727197, 25'd436318, -25'd2108872, 25'd1054436, 25'd181799, 25'd3381467, 25'd0}}, '{'{-25'd1599834, -25'd4472262, 25'd2945148, 25'd2726989, 25'd72720, -25'd3163308, -25'd690837, 25'd3272387, 25'd1490754}, '{25'd2545190, 25'd1527114, -25'd1636194, -25'd1599834, 25'd4363183, -25'd3017868, -25'd2472470, 25'd2981508, -25'd2908789}, '{-25'd2763349, -25'd981716, -25'd4181384, 25'd2108872, -25'd2690629, -25'd2981508, 25'd4145024, 25'd363599, 25'd2763349}, '{-25'd2690629, 25'd399958, 25'd2108872, 25'd1527114, 25'd2836069, -25'd2363391, 25'd3999584, 25'd1345315, 25'd727197}, '{25'd3999584, -25'd1599834, -25'd72720, -25'd4399543, -25'd1745273, 25'd3454186, 25'd4254103, 25'd3090588, -25'd1236235}, '{-25'd399958, 25'd1090796, 25'd2108872, -25'd2545190, -25'd981716, 25'd4035944, -25'd3526906, 25'd2181591, 25'd4363183}, '{-25'd1817993, 25'd145439, -25'd4654062, -25'd4544982, 25'd1854353, -25'd1599834, 25'd4035944, 25'd3708705, -25'd618118}, '{-25'd3526906, -25'd945356, -25'd4181384, 25'd872637, 25'd1672553, -25'd1563474, 25'd4472262, -25'd3126948, 25'd327239}, '{-25'd618118, -25'd36360, 25'd2581550, -25'd2799709, -25'd2581550, -25'd2072512, -25'd1345315, 25'd4617702, -25'd763557}}},
    '{'{'{25'd1852006, 25'd1997262, -25'd3885582, 25'd1634123, -25'd3050364, -25'd4030838, -25'd1270985, 25'd2723539, -25'd2687225}, '{25'd1525182, 25'd3268247, -25'd3994524, -25'd3014050, 25'd1053102, -25'd2142517, -25'd4176093, 25'd1852006, -25'd1852006}, '{25'd326825, 25'd2287773, 25'd835219, -25'd2433028, -25'd2106203, -25'd2142517, 25'd3086677, -25'd2433028, -25'd3921896}, '{25'd1234671, 25'd1561496, -25'd2106203, -25'd217883, 25'd2033576, -25'd1307299, 25'd1852006, -25'd1779379, 25'd4212407}, '{25'd581022, -25'd2360400, -25'd4430290, -25'd2469342, 25'd472080, 25'd3486130, -25'd835219, 25'd2578283, -25'd3740327}, '{-25'd2142517, 25'd2759853, 25'd3885582, -25'd2433028, 25'd3449816, 25'd1343613, 25'd1452554, 25'd3195619, 25'd1670437}, '{25'd3122991, 25'd2396714, -25'd4321348, -25'd3340874, -25'd1852006, -25'd1634123, 25'd3268247, -25'd2215145, -25'd1525182}, '{25'd3631385, 25'd2142517, 25'd3268247, 25'd835219, 25'd2033576, 25'd1053102, 25'd2505656, -25'd907846, -25'd4575545}, '{25'd2905108, 25'd2469342, -25'd2215145, -25'd726277, 25'd1307299, 25'd2796167, 25'd1852006, -25'd2215145, -25'd3122991}}, '{'{-25'd4248721, -25'd326825, 25'd2977736, -25'd798905, 25'd3486130, 25'd1198357, -25'd871532, 25'd4212407, 25'd1597809}, '{25'd581022, -25'd1452554, 25'd3921896, 25'd1307299, -25'd2505656, 25'd3449816, 25'd1125729, 25'd1053102, 25'd980474}, '{-25'd4067151, 25'd581022, 25'd2287773, -25'd2433028, 25'd3231933, -25'd4285035, 25'd1162043, -25'd2650911, -25'd3340874}, '{-25'd544708, -25'd3086677, 25'd1815693, 25'd2178831, -25'd798905, 25'd726277, 25'd1743065, -25'd3122991, -25'd1960948}, '{-25'd1053102, 25'd689963, -25'd1416240, 25'd544708, 25'd2868794, 25'd472080, 25'd3122991, 25'd3122991, -25'd290511}, '{25'd4176093, -25'd3994524, 25'd4139779, -25'd4176093, -25'd581022, -25'd1452554, 25'd2541970, -25'd2687225, 25'd3631385}, '{-25'd1234671, 25'd3014050, -25'd2541970, -25'd1053102, 25'd980474, 25'd1452554, -25'd3268247, 25'd689963, 25'd145255}, '{25'd2215145, 25'd508394, 25'd326825, 25'd1743065, -25'd1597809, 25'd0, 25'd3704013, -25'd653649, 25'd3449816}, '{25'd2469342, -25'd3377188, -25'd2941422, -25'd4176093, -25'd3449816, -25'd2977736, 25'd1779379, -25'd2215145, 25'd3159305}}, '{'{25'd1416240, 25'd1125729, 25'd980474, 25'd4611859, 25'd3122991, -25'd3086677, -25'd2178831, 25'd1924634, -25'd36314}, '{25'd3921896, 25'd4357662, 25'd4248721, -25'd1016788, -25'd2868794, 25'd72628, -25'd2905108, 25'd1234671, -25'd72628}, '{25'd3340874, -25'd3812954, -25'd1379926, -25'd1706751, -25'd2578283, -25'd472080, -25'd1416240, -25'd1343613, 25'd3776641}, '{-25'd2069890, 25'd2142517, 25'd2977736, -25'd145255, -25'd3014050, 25'd363139, -25'd4176093, 25'd4575545, -25'd108942}, '{-25'd145255, -25'd1561496, -25'd2977736, -25'd4648173, -25'd3522444, -25'd1561496, -25'd3885582, -25'd3413502, -25'd798905}, '{-25'd181569, -25'd2106203, -25'd4285035, -25'd3231933, -25'd3595071, -25'd1561496, 25'd435766, -25'd3667699, -25'd1089416}, '{25'd4067151, 25'd1198357, -25'd980474, -25'd3122991, -25'd1125729, 25'd3812954, 25'd399452, 25'd3667699, 25'd3704013}, '{-25'd2178831, 25'd0, 25'd3849268, 25'd1852006, -25'd4212407, -25'd472080, 25'd4176093, 25'd145255, -25'd2287773}, '{25'd871532, 25'd2142517, 25'd871532, -25'd3122991, -25'd653649, 25'd871532, 25'd2614597, 25'd1234671, 25'd4321348}}},
    '{'{'{25'd644620, 25'd2123456, -25'd4588181, 25'd2805995, 25'd606702, -25'd3981479, -25'd2426806, -25'd455026, 25'd1289241}, '{25'd75838, -25'd4853613, -25'd2047618, 25'd1971780, 25'd1023809, -25'd4588181, -25'd4133155, -25'd113757, -25'd2805995}, '{25'd1478835, 25'd1592592, 25'd3526453, -25'd1327160, -25'd1592592, -25'd113757, -25'd1365079, 25'd3829804, -25'd2047618}, '{25'd910052, -25'd3336859, 25'd1971780, 25'd3526453, 25'd3374778, -25'd758377, -25'd3336859, -25'd1706348, -25'd2388888}, '{-25'd4246911, -25'd3033508, -25'd1061728, 25'd3412697, 25'd2843914, -25'd4853613, 25'd758377, 25'd3261021, -25'd75838}, '{-25'd1213403, -25'd4019398, -25'd1630511, 25'd3147265, -25'd4360668, -25'd3678129, 25'd1365079, -25'd4588181, -25'd492945}, '{-25'd3336859, -25'd2805995, -25'd1023809, 25'd644620, -25'd151675, -25'd1251322, 25'd1251322, -25'd985890, -25'd3753966}, '{25'd2388888, 25'd2009699, 25'd2616401, -25'd4171074, 25'd1213403, -25'd3033508, -25'd2199293, 25'd113757, -25'd3185183}, '{-25'd341270, 25'd606702, 25'd151675, 25'd75838, 25'd303351, -25'd2047618, -25'd1251322, 25'd3261021, 25'd455026}}, '{'{-25'd568783, -25'd1744267, 25'd2843914, -25'd75838, 25'd4133155, 25'd265432, 25'd2692238, -25'd4853613, 25'd1440916}, '{25'd2843914, -25'd492945, 25'd1061728, 25'd189594, -25'd227513, -25'd341270, -25'd3298940, -25'd1820105, 25'd644620}, '{-25'd872134, -25'd3109346, -25'd3981479, 25'd3829804, -25'd758377, 25'd265432, -25'd4322749, 25'd872134, -25'd2388888}, '{25'd720458, 25'd3033508, 25'd4246911, 25'd189594, 25'd3147265, 25'd151675, -25'd2768076, -25'd455026, -25'd1554673}, '{-25'd2502644, 25'd4360668, -25'd2578482, -25'd3791885, -25'd1706348, -25'd720458, 25'd682539, -25'd3678129, -25'd1858024}, '{25'd2085537, 25'd189594, 25'd3791885, 25'd3109346, -25'd4095236, 25'd4474424, -25'd1971780, 25'd758377, -25'd2768076}, '{-25'd4133155, -25'd227513, 25'd1327160, -25'd1478835, 25'd379189, 25'd1137566, -25'd834215, -25'd2578482, -25'd2009699}, '{25'd3185183, 25'd872134, -25'd3526453, 25'd2464725, 25'd4095236, 25'd4133155, -25'd4853613, 25'd3147265, -25'd1630511}, '{-25'd1706348, 25'd1061728, 25'd0, -25'd3791885, 25'd910052, 25'd2843914, -25'd834215, 25'd2047618, -25'd3678129}}, '{'{-25'd492945, 25'd1933861, 25'd1213403, 25'd3943560, 25'd3109346, 25'd1744267, -25'd2881833, 25'd3223102, -25'd379189}, '{25'd530864, -25'd2881833, -25'd3905642, -25'd2881833, 25'd1289241, -25'd3716047, 25'd1630511, -25'd4853613, -25'd2085537}, '{25'd2540563, -25'd3298940, -25'd1061728, 25'd568783, -25'd2275131, 25'd1175484, 25'd1402997, 25'd3223102, 25'd2502644}, '{25'd3981479, -25'd227513, -25'd1592592, 25'd872134, -25'd2388888, 25'd4550262, -25'd4057317, -25'd2426806, 25'd2957670}, '{25'd265432, 25'd758377, 25'd3867723, 25'd3450615, -25'd3602291, -25'd3981479, 25'd2957670, 25'd910052, 25'd2995589}, '{-25'd1554673, -25'd3981479, 25'd4436506, 25'd151675, -25'd682539, -25'd1099647, -25'd2199293, -25'd4664019, -25'd985890}, '{-25'd872134, 25'd2009699, 25'd4246911, 25'd530864, 25'd265432, 25'd3374778, 25'd227513, -25'd3753966, -25'd3640210}, '{-25'd3716047, 25'd492945, 25'd2047618, 25'd4019398, 25'd341270, 25'd1099647, 25'd2578482, -25'd758377, 25'd1289241}, '{-25'd113757, -25'd4322749, 25'd2616401, -25'd3298940, 25'd2692238, -25'd2388888, -25'd417107, -25'd4436506, 25'd3336859}}},
    '{'{'{25'd593798, 25'd1543875, 25'd950077, -25'd2434572, -25'd237519, -25'd1425115, 25'd1068836, -25'd4572245, 25'd1068836}, '{-25'd4453485, 25'd3444028, 25'd59380, -25'd1603255, 25'd118760, 25'd3147129, 25'd1365735, 25'd415659, 25'd534418}, '{25'd534418, 25'd118760, -25'd178139, -25'd1959533, -25'd118760, 25'd415659, 25'd475038, -25'd2968990, -25'd1365735}, '{25'd2078293, 25'd2315812, -25'd2137673, 25'd2612711, 25'd712558, -25'd3978447, -25'd3919067, 25'd3147129, -25'd3622168}, '{25'd5344182, -25'd1781394, 25'd5047283, 25'd4750384, 25'd3622168, -25'd2553331, 25'd2553331, 25'd178139, -25'd1722014}, '{25'd950077, 25'd5106663, -25'd1306356, -25'd3800307, 25'd950077, -25'd3859687, 25'd2612711, -25'd3978447, -25'd1603255}, '{25'd2315812, 25'd1128216, -25'd2434572, -25'd2315812, -25'd3325269, -25'd4512865, -25'd3147129, 25'd356279, -25'd2078293}, '{25'd0, 25'd4037826, 25'd1009457, -25'd3740927, -25'd1603255, 25'd1068836, -25'd2850230, -25'd2137673, 25'd5225422}, '{25'd1009457, 25'd3919067, -25'd3265889, 25'd1603255, -25'd3681548, 25'd3740927, -25'd1543875, -25'd118760, 25'd4750384}}, '{'{-25'd1246976, 25'd2790851, -25'd534418, 25'd2078293, -25'd3800307, -25'd1009457, -25'd237519, 25'd2731471, -25'd4394105}, '{-25'd2731471, 25'd4750384, 25'd1543875, 25'd712558, 25'd2375192, 25'd3681548, -25'd1781394, -25'd4037826, -25'd2197053}, '{-25'd2790851, -25'd2078293, -25'd890697, -25'd1306356, -25'd3800307, -25'd4334725, 25'd4215966, -25'd1722014, 25'd1662634}, '{25'd831317, -25'd118760, 25'd2553331, 25'd3147129, -25'd4156586, -25'd2197053, 25'd1484495, -25'd3681548, -25'd3740927}, '{-25'd2612711, 25'd3740927, 25'd2553331, -25'd2493952, -25'd653178, 25'd2197053, -25'd3800307, 25'd1128216, 25'd2850230}, '{25'd4512865, 25'd1603255, -25'd593798, 25'd2018913, 25'd3147129, -25'd1840774, 25'd3978447, -25'd2315812, 25'd3206509}, '{-25'd1662634, -25'd2256432, -25'd4097206, -25'd1425115, -25'd7481855, -25'd3978447, 25'd4691004, 25'd475038, 25'd1543875}, '{25'd2137673, 25'd1306356, -25'd831317, 25'd1425115, -25'd5166043, 25'd1662634, -25'd534418, 25'd1365735, 25'd2375192}, '{25'd712558, 25'd2553331, -25'd2612711, 25'd59380, 25'd4215966, 25'd4631624, 25'd4453485, 25'd4512865, 25'd4037826}}, '{'{-25'd712558, 25'd2375192, 25'd1781394, 25'd4453485, -25'd3503408, -25'd2078293, 25'd1781394, 25'd2137673, 25'd4275346}, '{25'd3206509, 25'd1187596, 25'd3740927, -25'd3503408, 25'd2790851, -25'd1009457, -25'd1722014, 25'd3978447, 25'd2493952}, '{25'd1365735, 25'd296899, 25'd3740927, -25'd2137673, -25'd3978447, 25'd2315812, -25'd653178, 25'd3147129, -25'd1900154}, '{25'd2078293, -25'd3622168, -25'd5106663, -25'd2731471, -25'd5047283, -25'd1425115, 25'd1068836, 25'd4512865, 25'd4631624}, '{-25'd3562788, -25'd4512865, -25'd237519, -25'd5581701, -25'd7600614, 25'd237519, -25'd3800307, 25'd3681548, 25'd2790851}, '{25'd831317, 25'd1246976, -25'd2434572, -25'd2197053, -25'd6413018, -25'd1068836, -25'd2256432, 25'd890697, 25'd4869144}, '{25'd415659, 25'd2612711, 25'd1306356, -25'd593798, -25'd4928523, -25'd5819220, -25'd1722014, 25'd2018913, 25'd1840774}, '{-25'd534418, -25'd1662634, -25'd950077, -25'd4097206, -25'd2078293, 25'd2256432, -25'd3503408, 25'd4394105, 25'd4037826}, '{-25'd2078293, 25'd415659, 25'd1900154, -25'd1603255, -25'd4037826, 25'd3562788, 25'd4453485, 25'd4453485, -25'd1068836}}},
    '{'{'{-25'd179426, 25'd4234463, 25'd4485660, -25'd1327755, -25'd2942593, 25'd1399526, 25'd3660299, 25'd681820, -25'd2583740}, '{25'd4342119, 25'd2081346, -25'd1435411, -25'd3552643, -25'd3875610, 25'd3086134, 25'd4342119, 25'd466509, 25'd3050249}, '{25'd4557431, 25'd1255985, 25'd4126807, 25'd2045461, -25'd3624413, 25'd4198578, -25'd1794264, 25'd2476084, 25'd143541}, '{25'd4413890, -25'd3911496, 25'd3839725, 25'd1937805, 25'd4162693, -25'd3552643, -25'd789476, 25'd2081346, -25'd2727281}, '{-25'd2763167, 25'd1650723, -25'd1004788, -25'd1220100, 25'd3624413, -25'd1184214, -25'd466509, -25'd3193790, 25'd2691396}, '{25'd1112444, -25'd3911496, -25'd430623, -25'd143541, 25'd2296658, -25'd3480872, -25'd574164, 25'd2583740, 25'd143541}, '{25'd4342119, 25'd1076558, 25'd2476084, 25'd2799052, -25'd251197, 25'd1973690, -25'd2153117, 25'd2691396, -25'd2799052}, '{-25'd2691396, 25'd1866035, -25'd2224887, 25'd2296658, 25'd3014364, -25'd2978478, 25'd4055037, -25'd107656, 25'd143541}, '{-25'd1291870, 25'd2368429, -25'd1471297, 25'd322968, 25'd2476084, 25'd1650723, 25'd71771, -25'd1255985, -25'd933017}}, '{'{25'd538279, 25'd1255985, 25'd1830149, -25'd2799052, 25'd4449775, 25'd1291870, 25'd2511970, 25'd753591, 25'd3875610}, '{-25'd1004788, -25'd3588528, 25'd287082, 25'd394738, -25'd2189002, 25'd4306234, 25'd4342119, 25'd1901920, -25'd1830149}, '{-25'd1076558, 25'd3229675, 25'd4234463, 25'd2547855, 25'd3983266, -25'd1901920, 25'd2834937, -25'd2440199, -25'd1578952}, '{-25'd933017, -25'd2153117, 25'd1507182, -25'd3301446, 25'd1076558, -25'd2260773, 25'd1614838, 25'd4019151, -25'd3732069}, '{25'd3732069, -25'd3409102, -25'd143541, 25'd610050, 25'd2081346, 25'd215312, 25'd645935, -25'd2691396, 25'd2799052}, '{-25'd2117232, 25'd933017, 25'd3157905, 25'd466509, -25'd502394, 25'd1471297, 25'd3696184, 25'd3337331, 25'd3696184}, '{-25'd1866035, -25'd2870822, 25'd3875610, 25'd1291870, 25'd2476084, 25'd3767954, -25'd3086134, -25'd717706, -25'd2763167}, '{-25'd825361, -25'd2978478, -25'd2870822, -25'd1507182, -25'd4019151, -25'd3947381, 25'd2799052, -25'd2978478, 25'd2583740}, '{25'd71771, 25'd502394, 25'd4557431, -25'd1722493, 25'd358853, 25'd610050, -25'd3086134, 25'd143541, -25'd2727281}}, '{'{-25'd287082, 25'd1471297, 25'd4162693, 25'd3337331, -25'd358853, -25'd2727281, 25'd107656, 25'd1363641, -25'd3157905}, '{-25'd2511970, -25'd753591, 25'd968903, -25'd1650723, -25'd3696184, -25'd3480872, 25'd1937805, -25'd3193790, 25'd2870822}, '{-25'd3014364, -25'd2368429, -25'd1937805, 25'd1148329, -25'd394738, -25'd2045461, 25'd1758379, -25'd1507182, -25'd287082}, '{-25'd2727281, 25'd1686608, -25'd3696184, 25'd1291870, -25'd1399526, 25'd3086134, -25'd3265561, -25'd3947381, 25'd71771}, '{25'd1291870, -25'd1040673, -25'd215312, -25'd1148329, 25'd2511970, 25'd1507182, 25'd3050249, -25'd933017, 25'd1471297}, '{25'd1937805, 25'd3086134, 25'd1901920, -25'd3624413, 25'd1255985, 25'd1973690, -25'd3444987, -25'd2404314, -25'd1148329}, '{-25'd3983266, 25'd3839725, 25'd1363641, 25'd1399526, 25'd3193790, -25'd3947381, -25'd4019151, -25'd394738, 25'd430623}, '{-25'd3480872, 25'd1507182, 25'd3911496, -25'd2763167, -25'd3911496, -25'd2368429, -25'd1866035, 25'd4449775, 25'd1614838}, '{25'd3122019, 25'd287082, -25'd3229675, 25'd4198578, -25'd2619625, 25'd1184214, 25'd3480872, 25'd2117232, -25'd2511970}}},
    '{'{'{-25'd2354630, 25'd975490, -25'd2993744, -25'd1379141, -25'd3834684, -25'd3464670, 25'd2892832, 25'd1076402, 25'd1480053}, '{25'd1311866, 25'd1210953, 25'd3700133, -25'd3262845, 25'd3397395, 25'd4137422, 25'd2522818, 25'd3195570, -25'd1648241}, '{25'd1547329, -25'd908215, 25'd4204697, 25'd874577, 25'd2018255, 25'd1244590, -25'd1782792, 25'd2051892, -25'd2085530}, '{25'd3363758, 25'd1917342, -25'd1278228, 25'd2859194, -25'd201825, -25'd3868321, -25'd3767409, 25'd1110040, 25'd975490}, '{-25'd3330120, 25'd370013, 25'd302738, 25'd773664, 25'd302738, -25'd1883704, 25'd1446416, -25'd3767409, -25'd773664}, '{-25'd470926, -25'd2522818, -25'd3969234, 25'd1042765, 25'd370013, -25'd2623731, 25'd2388268, 25'd3027382, 25'd3700133}, '{25'd2320993, -25'd908215, 25'd168188, 25'd4070147, 25'd2724644, -25'd4070147, 25'd1345503, -25'd1446416, 25'd3632858}, '{-25'd1917342, -25'd2455543, 25'd235463, 25'd4137422, 25'd1984617, -25'd3969234, 25'd1244590, 25'd874577, 25'd605476}, '{-25'd908215, -25'd2623731, -25'd2186443, -25'd4238335, 25'd2926469, -25'd2287355, -25'd740027, -25'd2085530, -25'd706389}}, '{'{-25'd3061020, 25'd134550, -25'd1379141, -25'd3229207, -25'd504564, -25'd1917342, 25'd706389, 25'd2926469, -25'd1009127}, '{-25'd504564, 25'd2724644, -25'd3128295, -25'd2825556, -25'd2791919, -25'd1311866, -25'd874577, 25'd3565583, -25'd1816429}, '{25'd0, 25'd336376, 25'd1345503, -25'd538201, -25'd2623731, 25'd2791919, 25'd2152805, -25'd2051892, -25'd1480053}, '{25'd1715516, -25'd1614604, 25'd3262845, -25'd3262845, -25'd908215, -25'd4103784, 25'd2791919, -25'd2590093, -25'd4171060}, '{-25'd3363758, -25'd67275, 25'd3094657, -25'd908215, -25'd370013, 25'd2892832, 25'd1850067, -25'd1446416, 25'd908215}, '{-25'd4137422, -25'd1480053, -25'd1782792, 25'd538201, 25'd3565583, -25'd2892832, -25'd3061020, 25'd4271972, 25'd3767409}, '{-25'd2455543, -25'd235463, 25'd2522818, 25'd2859194, 25'd2489181, 25'd3128295, 25'd134550, 25'd538201, -25'd2489181}, '{-25'd2489181, 25'd2018255, 25'd571839, 25'd672752, -25'd1547329, 25'd4137422, 25'd2791919, -25'd874577, -25'd3969234}, '{-25'd3498308, 25'd3262845, -25'd1143678, -25'd2590093, -25'd168188, 25'd874577, -25'd3565583, 25'd33638, 25'd3195570}}, '{'{-25'd1950979, 25'd4070147, 25'd2657369, 25'd168188, 25'd3531946, -25'd3666496, -25'd2455543, -25'd3363758, 25'd100913}, '{-25'd2791919, 25'd3397395, 25'd2421906, 25'd3498308, 25'd1984617, 25'd2085530, 25'd1614604, 25'd1850067, 25'd1210953}, '{25'd370013, 25'd1311866, -25'd1412778, 25'd908215, 25'd269101, 25'd4238335, 25'd134550, 25'd3027382, 25'd3363758}, '{-25'd3901959, 25'd3363758, 25'd4036509, -25'd3397395, -25'd1782792, -25'd302738, 25'd302738, 25'd168188, 25'd941852}, '{25'd2825556, 25'd3801046, -25'd2522818, 25'd4070147, 25'd1749154, 25'd1177315, 25'd1850067, 25'd3262845, -25'd1547329}, '{25'd201825, 25'd2085530, -25'd3531946, 25'd4171060, 25'd3767409, -25'd2287355, 25'd3397395, -25'd4204697, 25'd1311866}, '{-25'd3901959, 25'd3262845, -25'd1076402, 25'd4238335, -25'd1950979, -25'd2993744, 25'd2993744, 25'd370013, -25'd235463}, '{-25'd3229207, 25'd1782792, 25'd2388268, 25'd3296483, 25'd2791919, -25'd201825, -25'd1816429, 25'd2455543, 25'd3161932}, '{-25'd1547329, 25'd3834684, 25'd1580966, -25'd1984617, 25'd2791919, 25'd672752, -25'd4204697, -25'd2691006, 25'd504564}}},
    '{'{'{25'd829725, -25'd2973182, -25'd3975767, -25'd3768336, 25'd3491760, 25'd898869, -25'd2973182, -25'd3768336, 25'd1002585}, '{25'd1970597, 25'd1348304, 25'd34572, -25'd3560904, -25'd691438, 25'd2385460, 25'd4390629, 25'd3699192, -25'd1313732}, '{25'd3664620, 25'd1071728, 25'd4183198, 25'd3872051, -25'd898869, 25'd864297, -25'd1763166, 25'd3630048, 25'd2212601}, '{25'd1624879, -25'd2696607, -25'd2938610, -25'd3076898, -25'd3007754, -25'd2938610, 25'd3249757, 25'd3664620, 25'd2212601}, '{-25'd1106300, -25'd2178029, -25'd2973182, 25'd1659450, 25'd829725, -25'd4079482, -25'd2765751, 25'd4321486, 25'd553150}, '{25'd2523748, -25'd1866882, 25'd4321486, -25'd172859, -25'd1140872, 25'd1728594, 25'd2178029, 25'd1037157, 25'd968013}, '{25'd691438, -25'd2350888, 25'd3699192, -25'd4010339, -25'd4010339, 25'd3837479, 25'd2316316, -25'd3249757, -25'd2385460}, '{25'd3664620, -25'd1348304, 25'd3215185, 25'd2178029, 25'd1244588, 25'd1486591, 25'd3422617, -25'd864297, -25'd518578}, '{-25'd414863, -25'd2938610, -25'd345719, 25'd2039741, 25'd3422617, -25'd4183198, 25'd138288, 25'd3906623, 25'd518578}}, '{'{25'd1313732, -25'd2869466, 25'd2385460, -25'd2523748, -25'd3872051, 25'd3768336, 25'd242003, -25'd484006, 25'd0}, '{-25'd1106300, -25'd3076898, -25'd3975767, 25'd760581, 25'd795153, -25'd242003, 25'd1486591, 25'd3664620, 25'd2834895}, '{-25'd3388045, 25'd2869466, 25'd2454604, -25'd1866882, 25'd3422617, 25'd4217770, -25'd1417447, 25'd3768336, 25'd345719}, '{-25'd2523748, -25'd1728594, 25'd829725, 25'd1417447, -25'd3111470, 25'd2039741, 25'd587722, -25'd311147, 25'd311147}, '{-25'd1140872, -25'd1348304, -25'd1071728, -25'd2592891, -25'd829725, 25'd1797738, 25'd3318901, 25'd2696607, -25'd2765751}, '{25'd172859, -25'd4114054, -25'd3422617, -25'd656866, -25'd3802907, -25'd1037157, -25'd1348304, 25'd172859, -25'd3699192}, '{25'd4010339, -25'd414863, -25'd3491760, 25'd3630048, 25'd4010339, -25'd1970597, -25'd553150, 25'd4010339, 25'd553150}, '{-25'd864297, 25'd4356058, 25'd1106300, 25'd345719, -25'd311147, 25'd4286914, 25'd2039741, 25'd4010339, -25'd138288}, '{25'd1348304, -25'd587722, -25'd2662035, 25'd553150, 25'd2592891, -25'd3664620, -25'd3491760, -25'd3975767, -25'd2350888}}, '{'{25'd311147, 25'd1659450, 25'd2800323, 25'd1244588, 25'd380291, -25'd2800323, -25'd4252342, -25'd3353473, 25'd4321486}, '{25'd726010, 25'd345719, 25'd3837479, 25'd587722, -25'd2869466, -25'd2005169, -25'd1071728, 25'd3630048, 25'd2039741}, '{-25'd1417447, -25'd484006, 25'd3215185, 25'd484006, 25'd311147, -25'd3630048, 25'd3284329, 25'd207431, 25'd2904038}, '{25'd2454604, -25'd2350888, 25'd4252342, -25'd3007754, -25'd2281744, 25'd1521163, 25'd3630048, -25'd4252342, 25'd2212601}, '{25'd4148626, -25'd3215185, -25'd1348304, 25'd3180613, -25'd2247173, 25'd1002585, 25'd3526332, 25'd2765751, -25'd1866882}, '{25'd1382875, -25'd933441, 25'd311147, -25'd829725, -25'd103716, 25'd1313732, -25'd1348304, -25'd3076898, 25'd3699192}, '{-25'd1175444, 25'd3422617, -25'd898869, 25'd3664620, 25'd3872051, 25'd1590307, -25'd2938610, -25'd2765751, 25'd4252342}, '{25'd726010, -25'd1624879, -25'd4010339, -25'd898869, 25'd3768336, 25'd3595476, 25'd4079482, 25'd1521163, 25'd3802907}, '{-25'd3180613, 25'd1486591, 25'd3560904, -25'd2627463, 25'd1037157, 25'd3007754, -25'd3802907, -25'd2592891, -25'd760581}}},
    '{'{'{-25'd4172177, 25'd4210454, -25'd1799012, 25'd1339690, -25'd2679380, 25'd2909041, -25'd4287008, -25'd2602826, 25'd995198}, '{25'd727260, 25'd1913843, -25'd76554, -25'd2373165, -25'd2832487, 25'd2717657, 25'd2487996, -25'd4057347, -25'd2296611}, '{25'd1799012, 25'd2526272, -25'd2909041, -25'd1913843, -25'd688983, -25'd2105227, -25'd2181781, 25'd1645905, 25'd1645905}, '{-25'd1454520, 25'd2296611, 25'd1186582, -25'd3636301, -25'd1760735, 25'd267938, 25'd4363561, 25'd3751132, 25'd306215}, '{25'd3100425, 25'd1339690, 25'd2641103, 25'd1799012, 25'd1684182, 25'd880368, 25'd267938, -25'd842091, 25'd1186582}, '{-25'd38277, 25'd688983, 25'd459322, 25'd4631499, 25'd2143504, 25'd1492797, -25'd1148306, -25'd1760735, 25'd2755933}, '{25'd3980793, 25'd3406640, 25'd1531074, 25'd1531074, 25'd3598024, -25'd76554, 25'd2487996, -25'd956921, -25'd2794210}, '{25'd2105227, 25'd727260, 25'd2755933, 25'd3942516, 25'd727260, 25'd3291809, 25'd4057347, 25'd4172177, -25'd2641103}, '{-25'd3827685, -25'd306215, 25'd1110029, 25'd4172177, -25'd2411442, 25'd535876, -25'd2641103, 25'd1722458, -25'd1416244}}, '{'{-25'd3980793, -25'd995198, -25'd2717657, -25'd918644, 25'd4401838, 25'd1148306, -25'd3559747, 25'd1033475, -25'd4172177}, '{25'd688983, -25'd3865962, 25'd2564549, -25'd4057347, -25'd2220058, 25'd3904239, -25'd4019070, -25'd2334888, 25'd2755933}, '{25'd1607628, -25'd1492797, 25'd2602826, -25'd688983, 25'd2487996, -25'd382769, 25'd1148306, 25'd2602826, -25'd2526272}, '{25'd1071752, 25'd1224859, 25'd1263136, 25'd4210454, 25'd4669776, -25'd2411442, -25'd1607628, -25'd2411442, -25'd1760735}, '{25'd2296611, 25'd3444917, 25'd4593222, 25'd3062148, 25'd612430, -25'd2641103, 25'd3521471, 25'd3827685, -25'd3138702}, '{25'd2947318, 25'd1837289, -25'd2947318, 25'd4861160, -25'd1454520, 25'd4478392, 25'd4133900, 25'd1607628, 25'd1952120}, '{-25'd842091, -25'd2947318, -25'd3559747, 25'd3712855, 25'd3406640, 25'd3674578, -25'd2296611, -25'd1263136, 25'd2296611}, '{-25'd1952120, -25'd2526272, -25'd2334888, 25'd2296611, 25'd114831, 25'd2181781, -25'd3674578, 25'd1377967, -25'd1186582}, '{-25'd2909041, -25'd918644, -25'd2105227, -25'd2449719, 25'd2487996, 25'd2258334, -25'd459322, 25'd3904239, -25'd956921}}, '{'{25'd3598024, 25'd2296611, 25'd1645905, -25'd3980793, 25'd267938, 25'd76554, 25'd2602826, 25'd2717657, 25'd114831}, '{25'd114831, 25'd1186582, 25'd2526272, -25'd2679380, 25'd497599, -25'd1263136, -25'd2909041, 25'd842091, -25'd1722458}, '{-25'd2679380, -25'd842091, 25'd2449719, 25'd2066950, 25'd2258334, -25'd2641103, -25'd4172177, 25'd1645905, -25'd2296611}, '{25'd4057347, 25'd650707, 25'd2870764, -25'd1990396, -25'd1531074, -25'd153107, -25'd3023871, 25'd995198, -25'd2794210}, '{-25'd2105227, 25'd76554, 25'd2028673, -25'd2641103, 25'd4095623, -25'd2181781, 25'd3904239, 25'd3942516, -25'd765537}, '{25'd3904239, 25'd382769, -25'd995198, -25'd1913843, 25'd382769, 25'd2985595, -25'd2143504, 25'd3215256, 25'd612430}, '{25'd1492797, 25'd956921, -25'd2487996, -25'd2641103, 25'd2296611, 25'd3980793, 25'd803814, -25'd2449719, 25'd3751132}, '{-25'd688983, 25'd4057347, -25'd1339690, 25'd4095623, 25'd2985595, 25'd1645905, -25'd76554, -25'd4401838, -25'd2870764}, '{-25'd3598024, -25'd1416244, -25'd1492797, 25'd956921, -25'd4287008, 25'd2641103, -25'd1875566, -25'd153107, 25'd2602826}}},
    '{'{'{-25'd804831, 25'd375588, 25'd804831, 25'd965797, -25'd2468148, 25'd3112012, 25'd1663317, 25'd4077809, -25'd2307182}, '{25'd1234074, 25'd965797, -25'd590209, 25'd2951046, 25'd375588, 25'd1126763, -25'd214622, -25'd590209, 25'd3863188}, '{25'd2199871, 25'd1609662, -25'd1019452, -25'd1180418, -25'd4882640, -25'd751175, -25'd4077809, -25'd3863188, 25'd4668018}, '{25'd1448695, -25'd2951046, 25'd1985249, -25'd1502351, 25'd1126763, -25'd1824283, 25'd3380289, -25'd697520, 25'd2360837}, '{-25'd3004702, -25'd3272978, -25'd2521803, -25'd2897391, -25'd4453397, -25'd1234074, -25'd5150917, 25'd214622, -25'd321932}, '{25'd1609662, -25'd912142, 25'd1770628, -25'd1073108, -25'd2629114, -25'd2360837, -25'd4131465, 25'd3648566, -25'd3433945}, '{25'd375588, -25'd1395040, -25'd2199871, 25'd643865, -25'd1716972, 25'd1931594, 25'd1985249, -25'd1234074, -25'd2468148}, '{-25'd536554, 25'd2951046, -25'd643865, 25'd1556006, -25'd643865, 25'd1287729, -25'd1931594, -25'd3809532, -25'd3326634}, '{25'd5419194, 25'd3648566, 25'd5902092, 25'd3594911, -25'd804831, 25'd3272978, 25'd6814234, -25'd160966, 25'd751175}}, '{'{-25'd1341385, -25'd1448695, 25'd2790080, -25'd4024154, 25'd1019452, 25'd1180418, 25'd3863188, -25'd1126763, -25'd3112012}, '{-25'd1019452, -25'd1341385, -25'd697520, -25'd2307182, 25'd4131465, -25'd2736425, 25'd2146215, 25'd3648566, -25'd1502351}, '{25'd536554, 25'd1073108, -25'd3165668, -25'd375588, -25'd643865, 25'd2038905, -25'd2575458, -25'd2253526, -25'd268277}, '{25'd53655, -25'd321932, -25'd1126763, 25'd268277, 25'd4077809, 25'd107311, 25'd3648566, -25'd1126763, -25'd53655}, '{-25'd3004702, 25'd2951046, -25'd2682769, -25'd5097262, -25'd2790080, -25'd590209, 25'd53655, 25'd751175, 25'd3702222}, '{-25'd2199871, -25'd2038905, 25'd4024154, 25'd2199871, 25'd2038905, 25'd965797, 25'd4453397, -25'd4507052, 25'd1609662}, '{25'd4721674, 25'd965797, 25'd2468148, 25'd268277, 25'd3326634, -25'd3272978, -25'd858486, -25'd3541255, 25'd3594911}, '{25'd4614363, -25'd4292431, -25'd4024154, -25'd5741126, 25'd4024154, 25'd160966, -25'd1770628, -25'd751175, 25'd2253526}, '{25'd4936295, 25'd3165668, -25'd3219323, 25'd1716972, 25'd697520, -25'd2575458, 25'd965797, -25'd3541255, -25'd2092560}}, '{'{25'd107311, 25'd160966, 25'd2521803, -25'd751175, -25'd2629114, -25'd2360837, 25'd536554, -25'd3970498, -25'd214622}, '{25'd1877938, 25'd2360837, -25'd482898, 25'd1931594, -25'd429243, -25'd2414492, -25'd1556006, 25'd1234074, -25'd590209}, '{-25'd2843735, 25'd2307182, -25'd321932, 25'd590209, -25'd268277, 25'd4399742, 25'd1824283, -25'd3916843, 25'd643865}, '{25'd160966, -25'd912142, 25'd3272978, -25'd912142, 25'd4024154, -25'd590209, 25'd3326634, -25'd2843735, 25'd2468148}, '{25'd160966, -25'd751175, -25'd1663317, 25'd4346086, 25'd1609662, 25'd2575458, 25'd5097262, -25'd2790080, -25'd804831}, '{-25'd1395040, 25'd3326634, 25'd1663317, 25'd3272978, 25'd3594911, 25'd1448695, 25'd3541255, 25'd2307182, -25'd1716972}, '{-25'd160966, -25'd4453397, -25'd107311, -25'd2951046, -25'd1877938, -25'd375588, 25'd429243, 25'd1770628, -25'd2360837}, '{-25'd4828985, -25'd1019452, -25'd3970498, -25'd107311, 25'd1395040, 25'd3058357, -25'd1019452, 25'd1985249, -25'd643865}, '{-25'd2575458, -25'd3594911, -25'd4989951, -25'd4292431, -25'd3004702, 25'd4346086, 25'd2897391, -25'd965797, -25'd2468148}}},
    '{'{'{-25'd2027841, -25'd2385696, 25'd2544742, 25'd397616, -25'd1351894, 25'd4373776, 25'd4254491, 25'd914517, -25'd3141166}, '{25'd3697828, -25'd516901, -25'd2902597, 25'd3538782, 25'd3220689, 25'd1749510, -25'd1232609, -25'd2743550, 25'd2107365}, '{-25'd1908557, 25'd1510941, 25'd3658067, 25'd2942358, -25'd1431417, 25'd3538782, 25'd914517, 25'd1510941, 25'd715709}, '{-25'd357854, 25'd4572584, -25'd1073563, 25'd4214729, -25'd159046, -25'd3777352, 25'd4015921, 25'd3141166, 25'd834994}, '{25'd1153086, 25'd3220689, -25'd1590464, 25'd3697828, 25'd3459259, -25'd79523, -25'd1232609, 25'd119285, -25'd357854}, '{-25'd3141166, 25'd1829033, 25'd4413537, -25'd3419497, -25'd477139, 25'd1272371, -25'd4373776, 25'd159046, -25'd3697828}, '{-25'd3141166, 25'd1630225, 25'd1988080, -25'd2823073, 25'd795232, -25'd3260451, -25'd4453299, -25'd4532822, -25'd3101405}, '{-25'd3936398, 25'd954278, -25'd2942358, 25'd1073563, 25'd994040, -25'd4095444, -25'd2465219, -25'd2544742, -25'd2027841}, '{25'd2902597, -25'd5089484, -25'd3697828, 25'd2703789, 25'd1908557, -25'd4334014, 25'd2385696, -25'd3976160, -25'd636186}}, '{'{-25'd4135206, -25'd2107365, -25'd3300213, 25'd397616, -25'd2783312, 25'd1590464, 25'd3419497, 25'd2743550, -25'd1391656}, '{25'd3379736, 25'd477139, -25'd2385696, -25'd1033802, 25'd397616, 25'd1033802, 25'd3220689, 25'd3180928, 25'd1948318}, '{25'd2664027, 25'd675947, 25'd3618305, 25'd4413537, 25'd4612345, -25'd914517, -25'd3419497, -25'd2902597, -25'd3817113}, '{-25'd3220689, -25'd3101405, 25'd2107365, 25'd2147126, 25'd2624265, -25'd3021881, 25'd1868795, 25'd4493060, 25'd2703789}, '{-25'd2306173, 25'd4055683, -25'd318093, -25'd39762, -25'd3618305, 25'd2902597, -25'd4453299, -25'd636186, 25'd4294252}, '{-25'd1312133, -25'd1550702, -25'd1391656, 25'd755470, -25'd2902597, 25'd556662, -25'd4055683, -25'd4135206, 25'd596424}, '{-25'd198808, 25'd1471179, 25'd2584504, 25'd3856875, -25'd1630225, -25'd1749510, -25'd3180928, 25'd3379736, -25'd2306173}, '{-25'd3180928, 25'd4214729, -25'd1113325, -25'd2544742, -25'd874755, 25'd3419497, -25'd3499020, 25'd2306173, 25'd2783312}, '{-25'd1988080, -25'd1192848, 25'd2544742, -25'd2107365, -25'd1829033, -25'd238570, 25'd2703789, -25'd357854, -25'd1550702}}, '{'{25'd3936398, 25'd477139, 25'd1192848, 25'd3658067, -25'd3061643, 25'd2266411, 25'd1351894, -25'd2942358, 25'd1630225}, '{25'd198808, 25'd2107365, -25'd1789272, 25'd1153086, -25'd1312133, 25'd596424, -25'd1391656, 25'd4493060, 25'd1391656}, '{-25'd2385696, -25'd4453299, -25'd3300213, -25'd1749510, -25'd755470, 25'd238570, 25'd3260451, 25'd2385696, -25'd1948318}, '{25'd2306173, -25'd1550702, -25'd4254491, -25'd3976160, -25'd1232609, -25'd119285, 25'd3697828, 25'd2982120, 25'd2743550}, '{25'd1988080, -25'd2504981, -25'd4453299, -25'd4691868, 25'd516901, -25'd954278, 25'd715709, -25'd3300213, -25'd2345934}, '{25'd1272371, 25'd3936398, 25'd2425457, 25'd1510941, 25'd2544742, -25'd3300213, 25'd3936398, 25'd516901, 25'd3936398}, '{-25'd1272371, 25'd3419497, 25'd1590464, -25'd2465219, -25'd4294252, 25'd1272371, -25'd4095444, 25'd715709, 25'd675947}, '{25'd3379736, 25'd357854, -25'd3379736, -25'd1272371, -25'd3379736, 25'd1312133, 25'd2862835, 25'd1829033, -25'd2823073}, '{25'd2266411, -25'd4015921, 25'd2186888, -25'd3737590, 25'd3856875, -25'd2664027, -25'd1073563, 25'd2743550, -25'd2504981}}},
    '{'{'{25'd4373227, 25'd2488828, -25'd2595493, -25'd3733243, 25'd3235477, 25'd2915485, 25'd1386633, 25'd1279969, -25'd3555469}, '{25'd1848844, 25'd2346610, -25'd2417719, -25'd391102, -25'd3733243, -25'd2631047, 25'd1955508, 25'd3235477, -25'd675539}, '{-25'd177773, -25'd3377696, 25'd1208860, 25'd2595493, -25'd3235477, 25'd71109, 25'd888867, -25'd2773266, 25'd4444337}, '{25'd639984, 25'd639984, 25'd2453274, -25'd3093258, 25'd3128813, 25'd4337672, 25'd2986594, 25'd2844375, -25'd2453274}, '{-25'd3911016, 25'd2559938, 25'd1564406, 25'd2453274, 25'd817758, 25'd3235477, 25'd1991063, 25'd3022149, -25'd3875461}, '{-25'd2239946, -25'd106664, -25'd1599961, 25'd4195454, -25'd3484360, 25'd2773266, -25'd2204391, -25'd3235477, 25'd924422}, '{25'd3306586, 25'd3128813, 25'd4408782, -25'd3128813, 25'd533320, 25'd2559938, 25'd319992, -25'd2986594, 25'd3057704}, '{25'd248883, -25'd1848844, -25'd3235477, 25'd2631047, -25'd319992, 25'd2417719, -25'd106664, -25'd817758, -25'd3022149}, '{25'd1599961, 25'd71109, 25'd1173305, 25'd2951039, -25'd3911016, 25'd1919953, 25'd3342141, 25'd2808821, -25'd3519915}}, '{'{-25'd959977, 25'd2879930, -25'd2631047, 25'd71109, -25'd2631047, -25'd3057704, -25'd2168836, 25'd2062172, 25'd782203}, '{25'd3377696, -25'd2702157, -25'd71109, 25'd675539, 25'd1137750, -25'd639984, 25'd3377696, 25'd2133282, -25'd995531}, '{-25'd3342141, -25'd782203, 25'd1422188, 25'd3484360, 25'd3591024, 25'd2559938, -25'd2915485, 25'd3484360, -25'd391102}, '{-25'd1671071, 25'd2773266, -25'd2773266, -25'd3519915, -25'd2773266, 25'd1919953, 25'd4515446, -25'd177773, -25'd3733243}, '{-25'd995531, 25'd2417719, 25'd2844375, -25'd675539, -25'd3875461, 25'd355547, 25'd4515446, 25'd4231008, -25'd1919953}, '{25'd2133282, -25'd2737711, 25'd2808821, 25'd1457742, -25'd3448805, -25'd2631047, -25'd319992, 25'd1066641, -25'd3022149}, '{-25'd142219, -25'd1137750, -25'd1884399, 25'd3804352, -25'd3164368, 25'd3804352, -25'd3164368, 25'd1386633, -25'd2453274}, '{-25'd746649, 25'd2488828, -25'd1244414, -25'd2524383, -25'd3377696, 25'd2275500, 25'd1813289, -25'd2062172, 25'd248883}, '{25'd3591024, 25'd2168836, -25'd782203, 25'd3982126, -25'd2311055, -25'd1457742, -25'd995531, -25'd319992, 25'd3093258}}, '{'{-25'd2133282, -25'd2879930, -25'd3982126, 25'd0, -25'd1102195, 25'd213328, 25'd1528852, -25'd2275500, -25'd3271032}, '{25'd3555469, -25'd3733243, 25'd0, 25'd2275500, 25'd3733243, -25'd319992, -25'd3235477, -25'd213328, -25'd2986594}, '{25'd3626579, -25'd2062172, 25'd2702157, -25'd2168836, -25'd853313, 25'd4231008, -25'd4088790, 25'd1137750, -25'd106664}, '{-25'd3235477, 25'd2488828, 25'd2026617, -25'd2453274, -25'd1031086, -25'd1457742, -25'd2417719, -25'd2239946, -25'd2737711}, '{-25'd3697688, 25'd106664, 25'd1137750, -25'd2239946, 25'd106664, 25'd2702157, -25'd3306586, 25'd3911016, -25'd675539}, '{25'd3768797, -25'd4088790, -25'd71109, 25'd2631047, -25'd1173305, -25'd248883, 25'd3911016, -25'd2773266, 25'd177773}, '{-25'd2488828, -25'd4017680, -25'd213328, -25'd2915485, -25'd1991063, 25'd0, 25'd1493297, 25'd3271032, -25'd1279969}, '{-25'd2275500, 25'd3199922, 25'd2702157, 25'd426656, -25'd462211, 25'd533320, 25'd2559938, 25'd1813289, 25'd1244414}, '{25'd3875461, 25'd4088790, 25'd1564406, 25'd4231008, 25'd2524383, -25'd3377696, -25'd462211, 25'd4515446, -25'd2844375}}},
    '{'{'{-25'd1729798, 25'd3036757, 25'd2075758, 25'd461279, 25'd3843996, 25'd1230079, -25'd4382155, -25'd38440, -25'd3228956}, '{25'd4228395, -25'd2229517, -25'd1960438, 25'd2267957, -25'd3498036, -25'd576599, 25'd538159, -25'd1499158, 25'd4189955}, '{-25'd461279, 25'd1960438, -25'd1729798, -25'd2652357, -25'd3344276, 25'd153760, 25'd4036195, -25'd2383277, -25'd1268519}, '{25'd3690236, -25'd307520, -25'd3767116, -25'd3651796, -25'd3267396, 25'd1537598, -25'd2652357, 25'd1537598, -25'd884119}, '{25'd1422278, 25'd4343715, 25'd2344837, -25'd3536476, 25'd1460718, -25'd1076319, -25'd1960438, 25'd153760, 25'd3574916}, '{25'd2075758, -25'd2767677, 25'd768799, -25'd1499158, -25'd3843996, 25'd4266835, 25'd1345398, -25'd2652357, -25'd3421156}, '{-25'd2344837, -25'd615039, 25'd1845118, -25'd192200, -25'd1076319, -25'd345960, 25'd2267957, 25'd768799, 25'd691919}, '{25'd4420595, 25'd3997755, 25'd2037318, -25'd230640, 25'd4382155, -25'd3690236, 25'd2037318, -25'd1614478, -25'd3228956}, '{-25'd76880, -25'd3305836, 25'd1921998, 25'd153760, -25'd2806117, -25'd1960438, 25'd884119, -25'd999439, -25'd2114198}}, '{'{-25'd1076319, -25'd2306397, 25'd3382716, 25'd2460157, -25'd461279, 25'd1499158, -25'd3574916, 25'd1191639, 25'd2959877}, '{25'd2690797, 25'd1306958, 25'd192200, 25'd1691358, -25'd2844557, 25'd2498597, 25'd1806678, 25'd2844557, -25'd2383277}, '{25'd1499158, -25'd3997755, -25'd1499158, -25'd2152638, -25'd2114198, -25'd2306397, -25'd3113636, 25'd2998317, 25'd2114198}, '{-25'd2767677, -25'd230640, 25'd4228395, -25'd3305836, -25'd2844557, -25'd2806117, -25'd115320, -25'd2882997, 25'd2075758}, '{-25'd269080, 25'd4266835, 25'd4420595, -25'd3613356, 25'd2921437, 25'd884119, -25'd2575477, 25'd2690797, 25'd653479}, '{25'd3152076, 25'd1806678, -25'd2191077, -25'd1768238, -25'd691919, -25'd2383277, 25'd884119, 25'd4113075, -25'd2690797}, '{25'd1652918, -25'd3190516, -25'd307520, -25'd3152076, -25'd1614478, 25'd3843996, 25'd2575477, -25'd922559, -25'd1537598}, '{-25'd2652357, -25'd269080, -25'd999439, -25'd3036757, -25'd2575477, 25'd76880, 25'd3728676, -25'd4382155, -25'd3228956}, '{25'd3574916, 25'd999439, 25'd115320, 25'd307520, 25'd2152638, -25'd1191639, 25'd192200, -25'd922559, 25'd4113075}}, '{'{-25'd1383838, 25'd2998317, -25'd2267957, 25'd2537037, -25'd2037318, 25'd1268519, -25'd3344276, 25'd1230079, -25'd2344837}, '{25'd3767116, -25'd807239, 25'd1460718, 25'd768799, -25'd1114759, -25'd1729798, -25'd3036757, -25'd3459596, 25'd922559}, '{-25'd38440, 25'd2537037, 25'd3113636, 25'd3882436, -25'd1883558, 25'd4535915, 25'd2959877, 25'd2267957, -25'd4036195}, '{-25'd1614478, -25'd3728676, -25'd1230079, 25'd4881874, -25'd1921998, 25'd3882436, 25'd4151515, -25'd115320, 25'd1499158}, '{25'd2229517, -25'd1960438, 25'd3728676, 25'd2152638, 25'd3228956, 25'd2191077, 25'd2498597, -25'd3882436, 25'd499719}, '{-25'd2729237, 25'd4343715, -25'd1576038, 25'd2537037, -25'd1845118, 25'd3613356, -25'd1921998, 25'd1921998, 25'd807239}, '{-25'd615039, -25'd768799, 25'd307520, -25'd2729237, 25'd4228395, 25'd3920875, 25'd2537037, -25'd2882997, 25'd1960438}, '{-25'd960999, -25'd2498597, 25'd3075196, 25'd1191639, 25'd4266835, 25'd768799, 25'd1806678, 25'd3613356, 25'd3113636}, '{-25'd1806678, -25'd3997755, 25'd1614478, 25'd3651796, 25'd4036195, 25'd538159, 25'd1691358, 25'd576599, 25'd307520}}},
    '{'{'{-25'd669319, -25'd739774, -25'd1303411, 25'd3346595, 25'd105682, 25'd3417050, -25'd2888640, 25'd2501139, 25'd176137}, '{25'd845456, -25'd3276140, -25'd2325003, -25'd246591, 25'd4403414, -25'd246591, 25'd3875005, 25'd2994322, 25'd1056819}, '{25'd2677276, 25'd669319, -25'd2642049, -25'd2007957, 25'd3910232, -25'd1514775, -25'd387500, -25'd1021592, -25'd4086368}, '{-25'd1021592, 25'd1197729, 25'd3804550, 25'd422728, -25'd1514775, 25'd3522731, 25'd880683, 25'd775001, 25'd3064776}, '{-25'd2148866, 25'd1127274, 25'd4438642, -25'd3381822, 25'd986365, -25'd1127274, 25'd3769323, -25'd3839777, 25'd3135231}, '{25'd4473869, -25'd880683, 25'd1796593, -25'd3593186, -25'd1268183, -25'd3240913, 25'd2888640, -25'd387500, -25'd2606821}, '{25'd70455, 25'd2888640, 25'd3769323, -25'd246591, -25'd1232956, 25'd2782958, -25'd3029549, -25'd563637, 25'd1796593}, '{-25'd704546, 25'd1479547, 25'd3135231, 25'd2571594, 25'd3734095, 25'd3417050, 25'd3276140, 25'd845456, -25'd1162501}, '{25'd915910, -25'd810228, -25'd3628413, 25'd1831820, -25'd3769323, 25'd2254548, 25'd1550002, 25'd1726138, 25'd1268183}}, '{'{25'd4086368, 25'd2642049, -25'd176137, 25'd0, -25'd634092, 25'd2642049, 25'd1162501, 25'd4438642, -25'd3417050}, '{-25'd3875005, 25'd1550002, -25'd2148866, 25'd4473869, -25'd1831820, -25'd2606821, 25'd2923867, -25'd1937502, -25'd1514775}, '{25'd1162501, 25'd4051141, 25'd2148866, -25'd3593186, 25'd1585229, -25'd2536367, 25'd669319, 25'd951137, -25'd3804550}, '{-25'd3839777, -25'd2536367, 25'd3311368, -25'd281819, 25'd246591, 25'd3205686, 25'd3064776, -25'd704546, 25'd1867048}, '{25'd3593186, 25'd3135231, 25'd1373865, 25'd1796593, -25'd4051141, 25'd493182, -25'd2325003, -25'd563637, -25'd775001}, '{-25'd3734095, -25'd4192050, 25'd3381822, -25'd1268183, 25'd1338638, 25'd1902275, 25'd3663641, -25'd3100004, -25'd669319}, '{-25'd2888640, 25'd3100004, -25'd387500, 25'd2007957, 25'd810228, 25'd3734095, -25'd3417050, 25'd1162501, -25'd246591}, '{-25'd3417050, 25'd3663641, 25'd457955, 25'd4262505, 25'd2677276, 25'd3029549, -25'd845456, -25'd2289775, 25'd4473869}, '{25'd3170458, 25'd739774, 25'd105682, -25'd528410, -25'd3910232, -25'd3734095, 25'd4332960, -25'd739774, -25'd3100004}}, '{'{-25'd2536367, 25'd3417050, 25'd493182, -25'd1514775, -25'd3417050, -25'd3100004, 25'd2501139, -25'd2007957, 25'd2325003}, '{-25'd3945459, -25'd2747731, 25'd211364, 25'd4403414, -25'd4262505, 25'd493182, 25'd1902275, -25'd3522731, 25'd3487504}, '{25'd3593186, 25'd3839777, -25'd2219321, 25'd317046, 25'd387500, 25'd2606821, 25'd3945459, -25'd2536367, -25'd2148866}, '{-25'd1127274, -25'd35227, 25'd3769323, -25'd4086368, -25'd3698868, -25'd281819, -25'd951137, -25'd1867048, -25'd2501139}, '{-25'd4368187, 25'd1092047, 25'd2078412, 25'd3452277, -25'd4227278, -25'd2818185, -25'd598864, -25'd3205686, 25'd3452277}, '{25'd3135231, 25'd2007957, 25'd3276140, -25'd1303411, 25'd1690911, -25'd2360230, -25'd2219321, 25'd775001, 25'd493182}, '{-25'd3593186, 25'd281819, 25'd3734095, -25'd2043184, -25'd2888640, 25'd951137, -25'd528410, 25'd352273, -25'd3346595}, '{25'd3804550, 25'd1127274, -25'd1162501, -25'd1444320, 25'd1444320, -25'd2747731, -25'd1690911, -25'd387500, 25'd3945459}, '{25'd493182, 25'd2606821, 25'd140909, -25'd1514775, -25'd1232956, -25'd810228, -25'd2219321, 25'd4368187, 25'd3135231}}},
    '{'{'{-25'd2480688, -25'd1386267, 25'd2407727, 25'd802576, 25'd1824036, 25'd1605151, 25'd4560089, -25'd1276825, -25'd839056}, '{25'd364807, -25'd4122320, 25'd4085840, 25'd839056, 25'd3830475, 25'd1094421, 25'd3246783, -25'd2918457, -25'd3684552}, '{-25'd1824036, 25'd1751074, -25'd839056, -25'd3246783, -25'd2334766, -25'd1787555, 25'd2042920, 25'd2444208, 25'd2225323}, '{25'd693134, -25'd2006439, 25'd4085840, 25'd3173822, 25'd1386267, -25'd1787555, -25'd1495709, -25'd1678113, 25'd2991418}, '{25'd2553650, 25'd2809015, -25'd1641632, -25'd1678113, -25'd1057941, -25'd2517169, -25'd1130902, -25'd2006439, -25'd729614}, '{-25'd2699573, 25'd3429187, 25'd4049359, 25'd3684552, -25'd3027899, -25'd1714593, -25'd3611590, 25'd3538629, 25'd4268243}, '{-25'd2699573, -25'd1313306, 25'd3173822, 25'd1386267, 25'd3392706, 25'd437769, 25'd3100861, 25'd1605151, -25'd766095}, '{25'd4122320, -25'd1969958, -25'd3392706, 25'd2371246, 25'd3246783, 25'd948499, -25'd547211, -25'd2918457, -25'd656653}, '{25'd547211, -25'd182404, -25'd656653, -25'd3939917, 25'd3137341, -25'd2663092, -25'd182404, 25'd2225323, -25'd547211}}, '{'{25'd1240344, 25'd4049359, 25'd1568671, 25'd875537, -25'd1751074, -25'd255365, -25'd3903436, 25'd693134, -25'd2553650}, '{-25'd3830475, 25'd802576, 25'd2225323, 25'd2663092, 25'd2480688, -25'd3027899, 25'd3575110, -25'd2809015, 25'd4085840}, '{-25'd1386267, 25'd2444208, -25'd1678113, 25'd3903436, -25'd2736053, 25'd1276825, 25'd255365, 25'd3137341, -25'd2371246}, '{-25'd1021460, 25'd2298285, -25'd3064380, -25'd3356225, 25'd4377685, 25'd1167383, -25'd2152362, 25'd4304724, -25'd437769}, '{-25'd948499, 25'd4231763, -25'd3429187, 25'd3976398, 25'd182404, 25'd2736053, 25'd4523608, 25'd4377685, -25'd839056}, '{-25'd3757513, -25'd2736053, 25'd1240344, 25'd2772534, -25'd1933478, 25'd474249, 25'd3173822, 25'd2845496, -25'd3903436}, '{25'd3210303, 25'd2188843, 25'd4268243, 25'd3283264, -25'd3538629, 25'd3429187, 25'd2480688, -25'd1824036, 25'd2079401}, '{25'd182404, -25'd510730, 25'd2772534, 25'd3611590, 25'd3684552, 25'd4633050, -25'd3976398, 25'd3793994, 25'd3721033}, '{-25'd1751074, -25'd510730, 25'd2954938, -25'd3721033, -25'd3538629, 25'd912018, 25'd4487128, -25'd3027899, 25'd3939917}}, '{'{-25'd2225323, -25'd1896997, -25'd2991418, 25'd3137341, -25'd3392706, 25'd948499, -25'd255365, 25'd984979, -25'd437769}, '{-25'd2407727, -25'd656653, -25'd2006439, 25'd182404, 25'd3465668, 25'd3173822, -25'd3684552, -25'd1240344, -25'd109442}, '{25'd3684552, -25'd2553650, 25'd4487128, 25'd2845496, -25'd620172, -25'd2444208, -25'd1787555, -25'd510730, -25'd3502148}, '{-25'd802576, 25'd3976398, 25'd255365, 25'd2225323, 25'd1641632, 25'd1276825, -25'd1094421, -25'd255365, 25'd328326}, '{25'd4523608, -25'd1240344, 25'd2772534, 25'd693134, 25'd1313306, -25'd109442, -25'd4158801, 25'd364807, -25'd3793994}, '{-25'd510730, 25'd218884, -25'd2553650, -25'd2772534, -25'd2371246, 25'd3793994, 25'd2261804, 25'd2006439, 25'd1021460}, '{25'd1203863, 25'd1459228, -25'd802576, -25'd3429187, -25'd72961, -25'd36481, 25'd3429187, -25'd364807, 25'd1678113}, '{25'd328326, -25'd2991418, -25'd4122320, 25'd2225323, 25'd2517169, -25'd547211, 25'd3137341, 25'd547211, 25'd4012878}, '{25'd802576, -25'd2444208, -25'd1860516, 25'd2115881, 25'd547211, -25'd2371246, 25'd2334766, -25'd2261804, 25'd3283264}}},
    '{'{'{25'd2166420, 25'd722140, -25'd1895618, 25'd4423108, 25'd2708025, 25'd90268, -25'd90268, -25'd2346955, 25'd1173478}, '{25'd0, 25'd2166420, 25'd90268, 25'd3520433, -25'd541605, -25'd2888560, 25'd992943, -25'd2346955, -25'd1805350}, '{-25'd1805350, -25'd2617758, 25'd4242573, 25'd6138191, 25'd1354013, -25'd6408993, -25'd1354013, 25'd3700968, -25'd2798293}, '{25'd4423108, -25'd270803, 25'd1173478, 25'd5686853, 25'd3700968, 25'd3159363, 25'd2076153, -25'd722140, 25'd451338}, '{25'd2708025, 25'd7311669, 25'd7131134, 25'd9207286, 25'd8936484, -25'd3069095, 25'd3881503, 25'd4423108, 25'd1354013}, '{-25'd6770063, -25'd1624815, -25'd1354013, 25'd4332841, 25'd1534548, -25'd2708025, -25'd7582471, -25'd2437223, -25'd8033809}, '{25'd1624815, 25'd270803, 25'd451338, 25'd3971771, 25'd992943, -25'd2346955, 25'd541605, -25'd5235516, -25'd180535}, '{-25'd1805350, 25'd631873, 25'd2888560, -25'd1173478, 25'd5506318, -25'd10471032, -25'd1715083, -25'd7401936, -25'd7763006}, '{-25'd180535, 25'd3700968, -25'd1715083, -25'd2617758, 25'd902675, -25'd11554242, -25'd4874446, -25'd2708025, -25'd1715083}}, '{'{-25'd4423108, -25'd3971771, -25'd3159363, -25'd180535, -25'd3159363, -25'd3700968, 25'd3791236, -25'd2888560, -25'd2798293}, '{25'd631873, 25'd2076153, 25'd1985885, -25'd4062038, 25'd361070, -25'd4693911, -25'd90268, 25'd4062038, -25'd3700968}, '{-25'd2076153, 25'd0, 25'd2076153, 25'd2076153, 25'd3159363, -25'd1083210, -25'd1173478, -25'd3430165, 25'd2166420}, '{-25'd2346955, -25'd1895618, 25'd1534548, -25'd2617758, 25'd5867388, -25'd3971771, 25'd2798293, 25'd3700968, 25'd2978828}, '{-25'd1083210, 25'd4062038, 25'd5506318, 25'd6860331, 25'd6318726, 25'd902675, 25'd4513376, 25'd1354013, -25'd1263745}, '{-25'd1624815, -25'd2708025, -25'd3881503, -25'd2256688, 25'd4152306, -25'd4152306, -25'd4513376, -25'd3610701, -25'd7311669}, '{-25'd3430165, -25'd4152306, -25'd1805350, -25'd2978828, -25'd992943, 25'd90268, 25'd2166420, -25'd3791236, -25'd3069095}, '{25'd1715083, 25'd1895618, 25'd180535, 25'd4513376, 25'd3520433, -25'd7040866, 25'd1895618, -25'd1715083, -25'd1715083}, '{-25'd2617758, -25'd4152306, 25'd3520433, -25'd722140, 25'd1263745, -25'd7131134, -25'd1263745, 25'd2617758, -25'd4603643}}, '{'{-25'd2798293, 25'd1173478, -25'd3159363, 25'd3430165, 25'd0, -25'd1083210, -25'd3069095, 25'd2256688, -25'd451338}, '{-25'd4332841, -25'd180535, -25'd1624815, 25'd2888560, 25'd1173478, -25'd1985885, -25'd2617758, -25'd1715083, 25'd3249630}, '{-25'd1895618, -25'd631873, -25'd2076153, -25'd2527490, 25'd2798293, -25'd992943, 25'd1805350, 25'd3159363, 25'd2888560}, '{25'd992943, 25'd90268, 25'd2527490, 25'd2527490, 25'd1985885, -25'd451338, 25'd4423108, 25'd5145248, 25'd1715083}, '{25'd5506318, 25'd180535, 25'd3339898, 25'd3430165, 25'd5596586, -25'd3069095, 25'd1173478, -25'd812408, 25'd180535}, '{-25'd5777121, -25'd1354013, 25'd722140, 25'd1173478, 25'd361070, -25'd5957656, -25'd4513376, -25'd5506318, -25'd6589528}, '{25'd992943, -25'd3249630, -25'd1263745, -25'd90268, 25'd2437223, -25'd5325783, -25'd2437223, 25'd2437223, 25'd1083210}, '{-25'd2888560, 25'd2708025, -25'd902675, 25'd4513376, 25'd4964713, -25'd4784178, 25'd2798293, -25'd4332841, 25'd90268}, '{-25'd2256688, 25'd3610701, 25'd2346955, -25'd1534548, -25'd541605, -25'd3610701, -25'd2437223, -25'd3700968, 25'd3069095}}},
    '{'{'{25'd2278134, -25'd1269780, -25'd4780347, 25'd2240787, 25'd3510567, 25'd1568551, -25'd3398528, 25'd2614252, -25'd3734646}, '{-25'd2875677, 25'd2950370, -25'd2502213, 25'd485504, 25'd4070764, -25'd4630961, 25'd1717937, -25'd3921378, -25'd1942016}, '{-25'd485504, 25'd2763638, -25'd3734646, 25'd336118, -25'd3884032, -25'd560197, -25'd3211795, 25'd1531205, -25'd336118}, '{25'd522850, -25'd3286488, -25'd149386, -25'd4780347, -25'd1045701, 25'd2352827, -25'd224079, 25'd2128748, -25'd2427520}, '{25'd3174449, -25'd2651598, 25'd2464866, 25'd1157740, -25'd672236, -25'd4182803, -25'd1008354, 25'd3547913, -25'd2166095}, '{25'd485504, 25'd37346, -25'd2091402, -25'd4481575, -25'd2091402, 25'd1456512, -25'd1867323, -25'd2763638, 25'd3361181}, '{-25'd3062410, -25'd149386, 25'd2576906, 25'd1568551, -25'd2838331, 25'd1942016, -25'd2950370, 25'd3622606, -25'd4145457}, '{25'd2278134, -25'd2838331, 25'd74693, 25'd896315, 25'd1307126, -25'd3697299, 25'd3697299, -25'd1829976, -25'd2464866}, '{25'd224079, -25'd1867323, -25'd4070764, -25'd1120394, -25'd3137102, 25'd1867323, -25'd4108110, 25'd3435874, 25'd2614252}}, '{'{-25'd4481575, -25'd3398528, 25'd1456512, -25'd1643244, 25'd3137102, -25'd3809339, 25'd2651598, -25'd4108110, 25'd1493858}, '{25'd373465, -25'd1717937, -25'd1269780, -25'd634890, 25'd2390173, -25'd1979362, 25'd3921378, -25'd3846685, -25'd149386}, '{-25'd1493858, -25'd2315480, -25'd2576906, -25'd896315, -25'd1867323, -25'd186732, 25'd373465, -25'd2502213, 25'd1867323}, '{25'd821622, -25'd1195087, -25'd4145457, -25'd3622606, -25'd3996071, 25'd1531205, 25'd3323835, 25'd2016709, 25'd3249142}, '{-25'd3286488, -25'd2987717, 25'd2128748, 25'd2240787, 25'd373465, 25'd3547913, -25'd3211795, -25'd2278134, 25'd3174449}, '{-25'd3025063, -25'd672236, -25'd1381819, 25'd1269780, 25'd410811, 25'd4257496, -25'd1307126, 25'd112039, 25'd1680591}, '{25'd4743000, 25'd2651598, -25'd2240787, 25'd1120394, -25'd2091402, 25'd1755284, 25'd1307126, -25'd2614252, 25'd560197}, '{-25'd3473221, 25'd2315480, 25'd1008354, -25'd2464866, 25'd1792630, 25'd2539559, -25'd1381819, 25'd3473221, 25'd1045701}, '{-25'd3249142, -25'd3846685, 25'd1792630, -25'd3435874, -25'd1867323, -25'd2054055, 25'd2016709, -25'd1120394, 25'd3025063}}, '{'{-25'd2614252, -25'd4780347, -25'd3734646, -25'd4406882, 25'd4182803, -25'd2166095, -25'd746929, -25'd522850, 25'd522850}, '{-25'd2464866, -25'd1120394, -25'd4182803, -25'd2950370, 25'd448157, -25'd2539559, 25'd224079, -25'd2464866, 25'd634890}, '{25'd3884032, -25'd634890, -25'd1232433, -25'd560197, 25'd186732, -25'd298772, -25'd4108110, 25'd2278134, -25'd1904669}, '{-25'd2502213, 25'd0, -25'd1531205, 25'd1605898, 25'd2278134, -25'd1643244, -25'd1045701, 25'd2427520, 25'd149386}, '{25'd4294843, -25'd3025063, 25'd3323835, 25'd1643244, 25'd112039, -25'd1456512, 25'd2427520, -25'd4033417, 25'd2315480}, '{25'd3884032, 25'd1269780, -25'd2278134, 25'd522850, -25'd261425, -25'd74693, -25'd1008354, 25'd1232433, 25'd3996071}, '{-25'd3510567, -25'd2800984, -25'd1120394, 25'd4518921, 25'd1456512, -25'd1045701, 25'd1717937, -25'd2054055, 25'd3547913}, '{25'd448157, 25'd4257496, 25'd2128748, 25'd2651598, 25'd1792630, 25'd4294843, 25'd4332189, -25'd1979362, -25'd485504}, '{-25'd560197, 25'd4257496, 25'd1419165, -25'd2203441, 25'd2240787, -25'd1419165, -25'd3921378, 25'd3062410, 25'd4145457}}},
    '{'{'{25'd1725667, 25'd4002079, -25'd1578802, -25'd2239696, 25'd2129547, 25'd2827157, -25'd2717008, 25'd1395220, 25'd3634916}, '{25'd1248355, 25'd844475, -25'd3671632, 25'd3745065, 25'd2276412, 25'd3010738, -25'd917908, -25'd1248355, -25'd3047455}, '{-25'd771043, -25'd1982681, 25'd954624, 25'd257014, 25'd734326, -25'd1285071, -25'd3377901, -25'd1174922, 25'd1872532}, '{-25'd146865, 25'd4332526, 25'd2863873, 25'd2019398, -25'd1799100, -25'd2239696, -25'd771043, 25'd4075511, 25'd624177}, '{-25'd807759, -25'd2092830, -25'd1652234, 25'd1578802, -25'd1285071, -25'd183582, 25'd3781781, 25'd3267752, -25'd3267752}, '{25'd550745, -25'd1505369, -25'd1872532, 25'd440596, -25'd3267752, -25'd4002079, 25'd1982681, -25'd1101490, 25'd991341}, '{-25'd771043, 25'd991341, -25'd3304469, -25'd440596, 25'd2459993, -25'd110149, -25'd4405958, 25'd330447, 25'd3708348}, '{-25'd3377901, 25'd2680291, -25'd146865, -25'd1762383, 25'd3671632, -25'd3451334, 25'd1064773, -25'd4699689, 25'd1542085}, '{-25'd514028, -25'd771043, 25'd440596, -25'd4479391, -25'd1982681, -25'd4259093, -25'd4479391, 25'd2423277, -25'd4479391}}, '{'{-25'd4002079, -25'd2092830, 25'd4112228, -25'd4222377, 25'd330447, -25'd2753724, -25'd4148944, 25'd2349844, 25'd1321788}, '{-25'd3524767, 25'd3598199, -25'd2496710, 25'd991341, 25'd4405958, -25'd3231036, -25'd1982681, 25'd3194320, -25'd3451334}, '{-25'd1285071, 25'd2386561, 25'd881192, 25'd477312, 25'd2900589, -25'd1138206, 25'd844475, 25'd403880, 25'd550745}, '{-25'd514028, 25'd2570142, 25'd477312, -25'd1835816, 25'd1395220, 25'd2680291, 25'd4148944, 25'd3341185, 25'd2533426}, '{-25'd4148944, 25'd2423277, -25'd3965363, -25'd2202979, -25'd3084171, -25'd2019398, 25'd3010738, -25'd4038795, -25'd1982681}, '{25'd844475, 25'd293731, -25'd2680291, 25'd330447, -25'd2386561, -25'd1688951, -25'd2533426, -25'd3194320, -25'd2386561}, '{-25'd183582, 25'd1945965, -25'd2570142, -25'd1578802, 25'd1945965, -25'd3010738, 25'd3267752, 25'd2790440, -25'd220298}, '{25'd1028057, -25'd954624, 25'd2459993, 25'd440596, 25'd917908, -25'd807759, 25'd2202979, 25'd2570142, 25'd2937306}, '{25'd2827157, -25'd3524767, -25'd917908, 25'd1028057, 25'd991341, -25'd550745, 25'd1725667, -25'd2937306, -25'd4699689}}, '{'{-25'd1652234, -25'd1285071, -25'd734326, 25'd4075511, 25'd3120887, 25'd2276412, 25'd2717008, 25'd1688951, 25'd734326}, '{25'd4038795, -25'd3855214, 25'd4112228, 25'd1174922, 25'd0, -25'd4038795, 25'd1762383, 25'd3634916, 25'd2753724}, '{-25'd3231036, 25'd4259093, 25'd3598199, -25'd1542085, -25'd3194320, -25'd1872532, -25'd3120887, -25'd4038795, -25'd1064773}, '{25'd4075511, -25'd2129547, 25'd3928646, 25'd2423277, 25'd1945965, -25'd3855214, 25'd3818497, 25'd2790440, 25'd330447}, '{25'd2423277, -25'd3708348, 25'd514028, 25'd36716, 25'd3891930, 25'd2056114, 25'd1578802, -25'd4112228, -25'd3377901}, '{-25'd1835816, -25'd771043, -25'd1909249, -25'd3524767, -25'd771043, 25'd2459993, 25'd1174922, 25'd2827157, 25'd3414618}, '{-25'd2056114, -25'd3084171, 25'd2166263, 25'd3781781, 25'd771043, -25'd514028, 25'd1615518, -25'd183582, 25'd1505369}, '{25'd3818497, 25'd1799100, 25'd1468653, 25'd1799100, 25'd3047455, -25'd2092830, 25'd1542085, -25'd697610, -25'd4699689}, '{-25'd4479391, 25'd1945965, -25'd4699689, -25'd4479391, -25'd3745065, -25'd2276412, -25'd1395220, -25'd1762383, -25'd3451334}}},
    '{'{'{-25'd246121, -25'd5845377, -25'd553773, -25'd1415196, -25'd4245589, 25'd1784378, -25'd2707332, -25'd1107545, -25'd3261105}, '{-25'd4860892, -25'd2215090, -25'd1230606, 25'd0, -25'd4430180, -25'd6091498, -25'd3999468, -25'd492242, -25'd4245589}, '{-25'd3445696, -25'd2584272, -25'd1722848, -25'd307651, -25'd5230074, -25'd3691817, -25'd7875876, -25'd7875876, 25'd123061}, '{25'd2215090, 25'd799894, -25'd861424, 25'd922954, -25'd4737832, -25'd4307120, -25'd5291604, -25'd5537725, 25'd61530}, '{-25'd3014984, 25'd3014984, -25'd2030499, -25'd123061, 25'd984484, -25'd3445696, -25'd2768863, 25'd430712, 25'd430712}, '{-25'd2338151, -25'd492242, -25'd2707332, -25'd4122529, -25'd4368650, -25'd984484, 25'd1784378, 25'd3630287, 25'd615303}, '{25'd1907439, -25'd4491711, 25'd1169075, 25'd492242, -25'd1907439, 25'd2461211, -25'd3753347, 25'd1353666, 25'd3199575}, '{-25'd3199575, -25'd4553241, 25'd3322635, -25'd984484, 25'd3814877, -25'd1046015, 25'd4368650, 25'd4553241, 25'd2030499}, '{25'd3568756, 25'd307651, 25'd1661318, -25'd2768863, -25'd1845908, 25'd123061, -25'd1784378, -25'd1907439, -25'd2645802}}, '{'{-25'd4368650, 25'd0, -25'd5353134, 25'd430712, -25'd369182, -25'd5045483, 25'd3568756, -25'd738363, 25'd3014984}, '{-25'd3445696, 25'd246121, -25'd2522742, -25'd3630287, -25'd5783846, 25'd1353666, -25'd2830393, -25'd5107013, -25'd1476727}, '{-25'd3507226, 25'd1538257, -25'd984484, 25'd3199575, -25'd3076514, -25'd1599787, -25'd4737832, 25'd738363, 25'd1107545}, '{-25'd1968969, -25'd1599787, 25'd369182, -25'd2584272, -25'd307651, 25'd2768863, 25'd4553241, -25'd3445696, 25'd3753347}, '{-25'd1230606, -25'd1661318, 25'd3261105, -25'd615303, 25'd0, 25'd4491711, 25'd4368650, 25'd307651, 25'd1169075}, '{-25'd492242, -25'd2707332, 25'd3691817, 25'd4860892, -25'd3384165, -25'd2399681, 25'd4184059, -25'd799894, 25'd4060999}, '{25'd1107545, 25'd1107545, 25'd3384165, 25'd2645802, 25'd1353666, 25'd3076514, 25'd4491711, 25'd2030499, 25'd2830393}, '{25'd4491711, 25'd4122529, 25'd4430180, 25'd3322635, -25'd1661318, 25'd5168544, 25'd738363, 25'd4553241, -25'd861424}, '{25'd3814877, 25'd676833, -25'd1353666, -25'd3014984, -25'd369182, 25'd5291604, 25'd1292136, 25'd1599787, -25'd676833}}, '{'{-25'd1845908, -25'd1415196, -25'd3691817, -25'd3014984, 25'd2399681, 25'd676833, -25'd3445696, 25'd984484, -25'd2891923}, '{-25'd2092030, -25'd3999468, -25'd1292136, -25'd5230074, -25'd7322103, -25'd6214558, -25'd7137513, -25'd6153028, -25'd6153028}, '{25'd2707332, -25'd3814877, 25'd2584272, -25'd2338151, 25'd799894, -25'd984484, -25'd246121, -25'd1538257, 25'd3199575}, '{25'd1169075, 25'd2215090, 25'd3568756, 25'd2645802, -25'd1476727, 25'd2645802, -25'd307651, 25'd4614771, -25'd2399681}, '{-25'd615303, 25'd615303, -25'd2338151, -25'd1476727, 25'd0, -25'd3138044, 25'd3014984, -25'd1722848, -25'd369182}, '{-25'd1415196, 25'd4060999, 25'd1599787, -25'd3568756, -25'd61530, 25'd3630287, 25'd3076514, 25'd799894, -25'd3691817}, '{-25'd3138044, 25'd1169075, -25'd1046015, -25'd4491711, -25'd2276620, 25'd2645802, -25'd3507226, 25'd1353666, 25'd4614771}, '{-25'd123061, 25'd369182, 25'd307651, 25'd2584272, 25'd123061, 25'd3507226, -25'd2461211, -25'd3568756, 25'd1230606}, '{-25'd2768863, -25'd922954, 25'd4368650, -25'd1169075, -25'd307651, -25'd3445696, -25'd2830393, 25'd3261105, 25'd984484}}},
    '{'{'{25'd2333639, -25'd382564, -25'd2983998, 25'd2792716, -25'd1185948, -25'd573846, -25'd1377230, 25'd2104101, 25'd2716203}, '{-25'd3519587, 25'd4322971, 25'd726871, -25'd2716203, -25'd3060510, 25'd573846, 25'd1759794, 25'd1568512, 25'd1989332}, '{-25'd3290049, 25'd3251792, -25'd3404818, 25'd1071179, 25'd3787382, -25'd459077, -25'd765128, 25'd3672613, 25'd879897}, '{-25'd1415486, -25'd1185948, -25'd1530255, 25'd3672613, -25'd497333, -25'd3557843, -25'd1759794, 25'd1338973, 25'd4208202}, '{25'd1989332, -25'd1453742, 25'd3519587, -25'd229538, 25'd1836306, 25'd1606768, 25'd2716203, -25'd994666, 25'd2907485}, '{25'd1491999, -25'd1798050, -25'd2524921, -25'd1606768, 25'd0, 25'd229538, 25'd0, -25'd3978664, -25'd420820}, '{-25'd3098767, -25'd2257126, 25'd2333639, 25'd2027588, 25'd4246458, 25'd2410152, 25'd4208202, 25'd229538, 25'd420820}, '{-25'd2448408, -25'd841640, 25'd1109435, -25'd191282, 25'd573846, 25'd3213536, 25'd2333639, 25'd994666, 25'd1606768}, '{-25'd38256, 25'd1071179, 25'd803384, 25'd573846, 25'd2486665, 25'd3902151, -25'd2677947, 25'd3710869, -25'd1912819}}, '{'{25'd4590766, 25'd3596100, -25'd3137023, 25'd382564, 25'd2180614, -25'd2639690, -25'd3863894, 25'd1415486, -25'd1645024}, '{25'd3557843, -25'd2716203, 25'd1530255, 25'd459077, 25'd2142357, 25'd956410, -25'd2869229, 25'd2104101, 25'd3672613}, '{-25'd2065845, 25'd306051, -25'd2371896, -25'd1683281, -25'd1300717, 25'd1338973, 25'd1721537, 25'd1491999, -25'd3787382}, '{25'd3137023, -25'd3902151, 25'd1836306, 25'd3213536, 25'd1147691, 25'd3863894, 25'd3060510, 25'd3710869, -25'd612102}, '{25'd612102, 25'd1568512, 25'd3902151, 25'd1683281, 25'd3672613, 25'd4284715, 25'd3825638, -25'd1147691, 25'd1530255}, '{-25'd726871, 25'd1109435, -25'd1759794, 25'd4858560, 25'd3443074, 25'd879897, -25'd1683281, 25'd573846, 25'd2716203}, '{25'd2869229, -25'd803384, 25'd344307, 25'd803384, 25'd1338973, -25'd3443074, -25'd1377230, -25'd1300717, -25'd3290049}, '{-25'd726871, -25'd2830972, -25'd3022254, 25'd1912819, 25'd2945741, -25'd3328305, 25'd1300717, 25'd2448408, -25'd1912819}, '{-25'd2601434, 25'd3710869, 25'd918153, 25'd459077, -25'd3902151, -25'd2677947, 25'd1109435, -25'd3557843, 25'd1491999}}, '{'{25'd1989332, 25'd4399484, -25'd2639690, 25'd4437740, -25'd1032922, -25'd650358, -25'd3710869, -25'd191282, 25'd3366561}, '{-25'd2792716, -25'd535589, -25'd2180614, -25'd3290049, 25'd2180614, -25'd1721537, -25'd3481331, -25'd879897, 25'd4093433}, '{25'd2524921, 25'd3443074, -25'd1109435, 25'd3863894, -25'd841640, 25'd3443074, 25'd420820, 25'd3940407, -25'd3557843}, '{-25'd1874563, -25'd2983998, 25'd1721537, 25'd2371896, -25'd3940407, -25'd2333639, 25'd688615, 25'd497333, -25'd3213536}, '{25'd535589, -25'd3366561, 25'd3902151, -25'd2333639, 25'd2677947, 25'd535589, -25'd3137023, 25'd3290049, 25'd765128}, '{25'd2601434, -25'd803384, 25'd1568512, 25'd1759794, -25'd191282, -25'd1300717, 25'd2218870, 25'd3213536, -25'd2907485}, '{-25'd2907485, 25'd1147691, 25'd3022254, -25'd535589, -25'd841640, -25'd535589, 25'd3863894, 25'd1338973, -25'd956410}, '{25'd229538, -25'd459077, -25'd573846, 25'd4361227, -25'd1224204, -25'd3098767, 25'd1645024, 25'd2869229, -25'd1224204}, '{-25'd2486665, 25'd3328305, -25'd3175280, -25'd1645024, -25'd2830972, -25'd2639690, 25'd2027588, 25'd994666, -25'd420820}}}
};
