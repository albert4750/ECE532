localparam bit signed [0:10][31:0] Bias = '{-32'd12125, -32'd20934, -32'd15439, 32'd29802, -32'd24375, 32'd23852, -32'd14579, 32'd15225, -32'd30906, 32'd8742, 32'd3751};
