localparam bit signed [0:10][15:0] Output8 = '{-16'd5612, -16'd20672, -16'd10219, -16'd11403, -16'd9779, 16'd24723, -16'd4279, 16'd17134, -16'd6047, -16'd4199, 16'd17051};
