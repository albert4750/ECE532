localparam bit signed [0:2][0:31][0:4][0:4][24:0] Weight3 = '{
    '{'{'{-25'd837, 25'd1883, 25'd2929, 25'd2302, 25'd4185}, '{25'd0, 25'd2720, 25'd2720, 25'd2511, -25'd418}, '{-25'd628, 25'd3139, 25'd837, 25'd2511, 25'd1674}, '{25'd3766, 25'd1674, 25'd209, 25'd0, 25'd1465}, '{25'd0, 25'd1255, 25'd2511, 25'd209, 25'd3348}}, '{'{25'd10671, 25'd7742, 25'd6905, 25'd5859, 25'd6696}, '{25'd7951, 25'd4813, 25'd6696, 25'd4813, 25'd6277}, '{25'd4603, 25'd5859, 25'd2302, 25'd5231, 25'd2092}, '{25'd3348, 25'd2929, 25'd1883, 25'd5650, 25'd6486}, '{25'd5859, 25'd3139, 25'd6068, 25'd5650, 25'd4603}}, '{'{-25'd1046, 25'd2511, 25'd2929, 25'd2929, 25'd2511}, '{25'd3348, 25'd3348, 25'd3348, 25'd2929, 25'd2720}, '{25'd0, 25'd1674, 25'd2511, 25'd1255, -25'd209}, '{25'd0, -25'd1046, 25'd1883, 25'd837, 25'd1255}, '{-25'd418, 25'd837, 25'd209, 25'd0, 25'd2929}}, '{'{25'd1883, 25'd2511, 25'd4603, 25'd2511, 25'd3976}, '{25'd5231, 25'd4185, 25'd1255, 25'd1465, 25'd1255}, '{25'd1674, 25'd5022, 25'd3557, 25'd2302, 25'd628}, '{25'd5022, 25'd2929, 25'd3139, 25'd2511, 25'd1465}, '{25'd1674, 25'd4185, 25'd3139, 25'd3766, 25'd3766}}, '{'{25'd5650, 25'd5022, 25'd4185, 25'd1465, 25'd5022}, '{25'd5022, 25'd4185, 25'd4813, 25'd3557, 25'd1674}, '{25'd5231, 25'd5650, 25'd4185, 25'd2302, 25'd5231}, '{25'd8579, 25'd3139, 25'd6486, 25'd3766, 25'd6905}, '{25'd8370, 25'd5859, 25'd4394, 25'd2302, 25'd3139}}, '{'{25'd4185, 25'd20924, 25'd26574, 25'd16321, 25'd14856}, '{-25'd2511, 25'd16739, 25'd20715, 25'd7742, 25'd9416}, '{25'd25946, 25'd26574, 25'd26574, 25'd25737, 25'd26574}, '{25'd7114, 25'd17576, 25'd18204, 25'd10881, 25'd12554}, '{-25'd2929, 25'd7951, 25'd9834, -25'd837, 25'd1883}}, '{'{-25'd418, -25'd1046, -25'd1046, 25'd1046, 25'd1255}, '{25'd1674, -25'd837, 25'd1674, 25'd1883, 25'd1465}, '{25'd418, 25'd418, -25'd209, -25'd628, 25'd2511}, '{25'd2720, 25'd628, -25'd418, -25'd837, 25'd0}, '{25'd628, 25'd1465, 25'd418, 25'd1046, 25'd1255}}, '{'{-25'd1255, -25'd3348, -25'd2511, -25'd209, -25'd3976}, '{-25'd418, -25'd4813, -25'd3766, -25'd4394, -25'd2092}, '{-25'd3348, -25'd4394, -25'd3766, -25'd418, -25'd1046}, '{-25'd837, -25'd2720, -25'd1465, -25'd418, -25'd209}, '{-25'd4185, -25'd3139, -25'd5022, -25'd1465, -25'd4603}}, '{'{-25'd1046, 25'd209, -25'd628, 25'd837, 25'd0}, '{-25'd418, 25'd1046, 25'd0, 25'd1465, 25'd3139}, '{25'd3348, 25'd1046, 25'd1883, -25'd1046, 25'd1883}, '{-25'd628, 25'd1465, 25'd2092, 25'd1465, 25'd209}, '{25'd1883, 25'd3139, 25'd3139, -25'd1255, 25'd209}}, '{'{25'd14019, 25'd10462, 25'd13182, 25'd12973, 25'd14228}, '{25'd15275, 25'd8788, 25'd10881, 25'd12554, 25'd13391}, '{25'd12554, 25'd10462, 25'd12345, 25'd13182, 25'd10881}, '{25'd11927, 25'd9625, 25'd8997, 25'd12973, 25'd14019}, '{25'd13810, 25'd7951, 25'd9207, 25'd13601, 25'd10671}}, '{'{25'd4185, 25'd1255, 25'd5022, 25'd4185, 25'd5859}, '{25'd4813, 25'd5022, 25'd3976, 25'd4394, 25'd5231}, '{25'd2511, 25'd1465, 25'd837, 25'd3557, 25'd4185}, '{25'd5231, 25'd3557, 25'd4185, 25'd1046, 25'd2511}, '{25'd3348, 25'd1046, 25'd2929, 25'd1046, 25'd5650}}, '{'{-25'd628, 25'd2302, 25'd0, 25'd3348, 25'd1255}, '{25'd3557, 25'd3766, 25'd1046, 25'd2511, 25'd1674}, '{25'd2302, -25'd628, 25'd3976, -25'd418, 25'd1674}, '{25'd3348, -25'd628, 25'd1674, 25'd1674, 25'd3766}, '{25'd3976, 25'd628, 25'd1046, 25'd1883, 25'd2720}}, '{'{25'd3557, 25'd6486, 25'd5859, 25'd5022, 25'd1674}, '{25'd3139, 25'd5231, 25'd2720, 25'd1255, 25'd4813}, '{25'd2720, 25'd2720, 25'd6068, 25'd3348, 25'd6486}, '{25'd4603, 25'd3976, 25'd3976, 25'd3976, 25'd5650}, '{25'd3557, 25'd4394, 25'd3976, 25'd3348, 25'd3139}}, '{'{25'd1255, 25'd3348, 25'd209, -25'd837, 25'd1883}, '{-25'd418, 25'd2720, -25'd1046, 25'd1046, 25'd3348}, '{25'd3557, 25'd1046, -25'd628, -25'd209, 25'd837}, '{-25'd1046, 25'd3139, 25'd837, 25'd1046, 25'd1883}, '{25'd2511, -25'd837, -25'd1046, -25'd418, 25'd0}}, '{'{25'd3348, 25'd3348, 25'd209, 25'd1883, 25'd0}, '{25'd837, 25'd1465, 25'd2092, -25'd628, 25'd2929}, '{-25'd209, 25'd2929, -25'd837, -25'd1465, 25'd2092}, '{25'd2511, 25'd837, 25'd837, 25'd209, 25'd1046}, '{-25'd418, 25'd837, 25'd2720, 25'd1883, -25'd418}}, '{'{25'd5859, 25'd5650, 25'd2720, 25'd3139, 25'd1465}, '{25'd6068, 25'd2720, 25'd1465, -25'd209, 25'd3766}, '{25'd7742, 25'd5231, 25'd2720, 25'd4185, 25'd418}, '{25'd3139, 25'd1046, 25'd628, -25'd209, 25'd3976}, '{25'd4603, 25'd2302, 25'd5859, 25'd6277, 25'd8370}}, '{'{25'd4394, 25'd3766, 25'd4394, 25'd3766, 25'd5859}, '{25'd5231, 25'd5022, 25'd4185, 25'd3348, 25'd3766}, '{25'd6696, 25'd3139, 25'd5022, 25'd6486, 25'd6486}, '{25'd7323, 25'd3348, 25'd6486, 25'd6277, 25'd4394}, '{25'd2929, 25'd5859, 25'd8160, 25'd7742, 25'd3976}}, '{'{25'd1883, 25'd5859, 25'd4813, 25'd4603, 25'd5440}, '{25'd5022, 25'd3766, 25'd3557, 25'd2929, 25'd7323}, '{25'd4813, 25'd4394, 25'd2511, 25'd4394, 25'd4394}, '{25'd4185, 25'd6068, 25'd3766, 25'd2302, 25'd2092}, '{25'd7114, 25'd6277, 25'd1465, 25'd1046, 25'd628}}, '{'{-25'd5231, -25'd628, -25'd3348, -25'd3557, -25'd2929}, '{-25'd4185, -25'd3976, -25'd4603, -25'd1255, -25'd2720}, '{-25'd2302, -25'd1046, -25'd3976, -25'd2511, -25'd1046}, '{-25'd2720, -25'd1255, -25'd2929, -25'd628, -25'd5650}, '{-25'd5022, -25'd418, -25'd3976, -25'd1883, -25'd5231}}, '{'{25'd22807, 25'd26364, 25'd25527, 25'd24272, 25'd20087}, '{25'd20715, 25'd23644, 25'd21133, 25'd19459, 25'd12554}, '{25'd16321, 25'd21133, 25'd16112, 25'd16739, 25'd11090}, '{25'd15902, 25'd13601, 25'd17367, 25'd16112, 25'd9625}, '{25'd18413, 25'd16949, 25'd18413, 25'd17158, 25'd12345}}, '{'{25'd11718, 25'd11299, 25'd12764, 25'd12764, 25'd13601}, '{25'd12554, 25'd10253, 25'd8997, 25'd12136, 25'd9416}, '{25'd11718, 25'd13182, 25'd9416, 25'd12764, 25'd10253}, '{25'd12136, 25'd12136, 25'd10671, 25'd8997, 25'd11299}, '{25'd15275, 25'd14019, 25'd10881, 25'd12345, 25'd9625}}, '{'{25'd209, 25'd1674, 25'd3976, 25'd3976, 25'd4813}, '{25'd2511, 25'd0, -25'd837, 25'd2929, 25'd3976}, '{25'd1046, 25'd628, 25'd2929, 25'd4185, 25'd2511}, '{25'd1046, -25'd1046, 25'd4185, 25'd1255, 25'd3348}, '{25'd3348, 25'd2720, 25'd4813, 25'd2720, 25'd6068}}, '{'{-25'd6905, -25'd418, 25'd2302, -25'd2511, -25'd1674}, '{25'd7533, 25'd15484, 25'd15484, 25'd17158, 25'd16530}, '{25'd15693, 25'd19459, 25'd23226, 25'd22180, 25'd26364}, '{25'd8160, 25'd14647, 25'd15693, 25'd15275, 25'd18832}, '{25'd5650, 25'd10671, 25'd12973, 25'd10671, 25'd20296}}, '{'{25'd8997, 25'd12764, 25'd10044, 25'd11508, 25'd12554}, '{25'd11508, 25'd10253, 25'd10881, 25'd11090, 25'd7323}, '{25'd7951, 25'd10253, 25'd9207, 25'd9416, 25'd10253}, '{25'd7323, 25'd11090, 25'd8997, 25'd11718, 25'd8160}, '{25'd9207, 25'd10253, 25'd9416, 25'd8370, 25'd11299}}, '{'{25'd4394, 25'd4813, 25'd4394, 25'd3976, 25'd6277}, '{25'd6068, 25'd4813, 25'd6696, 25'd5440, 25'd5650}, '{25'd7742, 25'd5440, 25'd8579, 25'd8997, 25'd12554}, '{25'd8579, 25'd8997, 25'd11299, 25'd7742, 25'd13391}, '{25'd12136, 25'd9834, 25'd11718, 25'd10253, 25'd14438}}, '{'{25'd10253, 25'd11718, 25'd12554, 25'd8997, 25'd12764}, '{25'd10253, 25'd10462, 25'd11718, 25'd9834, 25'd9416}, '{25'd10671, 25'd11299, 25'd8788, 25'd10881, 25'd13391}, '{25'd12554, 25'd11927, 25'd9834, 25'd9834, 25'd11299}, '{25'd15275, 25'd12345, 25'd12136, 25'd11927, 25'd10671}}, '{'{25'd11508, 25'd8788, 25'd8997, 25'd8579, 25'd12764}, '{25'd11508, 25'd11299, 25'd11927, 25'd7951, 25'd9834}, '{25'd8788, 25'd10462, 25'd11090, 25'd9416, 25'd9625}, '{25'd10671, 25'd12345, 25'd11508, 25'd7323, 25'd8370}, '{25'd10671, 25'd10253, 25'd7951, 25'd8788, 25'd8160}}, '{'{25'd2092, 25'd1255, 25'd3139, -25'd209, 25'd1465}, '{25'd3976, 25'd418, 25'd628, 25'd3557, 25'd2092}, '{25'd0, 25'd418, 25'd1465, 25'd1255, 25'd1255}, '{25'd3348, 25'd1255, 25'd628, 25'd1255, 25'd4813}, '{25'd0, 25'd3766, 25'd4603, 25'd2720, 25'd1674}}, '{'{25'd5650, 25'd5022, 25'd3348, 25'd2092, 25'd4185}, '{25'd2511, 25'd3557, 25'd3348, 25'd4813, 25'd6486}, '{25'd1255, 25'd4813, 25'd5231, 25'd4185, 25'd7323}, '{25'd3766, 25'd4603, 25'd2511, 25'd7742, 25'd6486}, '{25'd2720, 25'd6277, 25'd5859, 25'd7951, 25'd6068}}, '{'{25'd1046, 25'd837, 25'd209, 25'd2302, 25'd3139}, '{-25'd418, 25'd1465, 25'd2929, 25'd2720, 25'd1465}, '{25'd2092, 25'd0, 25'd837, -25'd418, 25'd2929}, '{25'd3557, 25'd209, 25'd2092, 25'd3766, 25'd209}, '{25'd1674, 25'd837, 25'd3348, 25'd1046, 25'd3766}}, '{'{25'd7323, 25'd5440, 25'd2929, 25'd1883, 25'd2302}, '{25'd6696, 25'd3976, 25'd2720, 25'd5231, 25'd2511}, '{25'd5231, 25'd3139, 25'd1255, 25'd628, 25'd5440}, '{25'd5859, 25'd4813, 25'd3976, 25'd1674, 25'd6277}, '{25'd7114, 25'd7114, 25'd3766, 25'd2302, 25'd6068}}, '{'{25'd12973, 25'd10671, 25'd15275, 25'd15275, 25'd17158}, '{25'd11508, 25'd8370, 25'd11090, 25'd14647, 25'd15065}, '{25'd11299, 25'd10881, 25'd9834, 25'd15484, 25'd16112}, '{25'd11508, 25'd8997, 25'd13182, 25'd15693, 25'd13601}, '{25'd12764, 25'd11090, 25'd14228, 25'd16530, 25'd15275}}},
    '{'{'{-25'd197, -25'd197, -25'd197, 25'd1577, 25'd3154}, '{-25'd197, 25'd394, 25'd3154, 25'd1183, 25'd3745}, '{25'd2366, -25'd394, 25'd3745, 25'd4140, 25'd394}, '{25'd0, 25'd591, 25'd2957, 25'd4140, 25'd2366}, '{25'd4534, 25'd2366, 25'd2760, 25'd3745, 25'd197}}, '{'{25'd9265, 25'd7294, 25'd6702, 25'd5322, 25'd4140}, '{25'd6111, 25'd2366, 25'd6505, 25'd2563, 25'd6900}, '{25'd6505, 25'd2957, 25'd2366, 25'd4337, 25'd4731}, '{25'd4140, 25'd4337, 25'd2168, 25'd2760, 25'd7688}, '{25'd4337, 25'd6308, 25'd3943, 25'd4731, 25'd8082}}, '{'{25'd197, 25'd3154, 25'd0, 25'd986, 25'd197}, '{-25'd986, 25'd1577, 25'd3351, 25'd3548, -25'd789}, '{25'd1380, 25'd1971, 25'd394, 25'd3154, 25'd3548}, '{25'd1183, -25'd789, -25'd197, 25'd1577, -25'd197}, '{-25'd789, 25'd197, 25'd0, 25'd0, 25'd2168}}, '{'{25'd986, 25'd394, 25'd4534, 25'd1774, 25'd1183}, '{25'd4337, 25'd1774, 25'd2760, 25'd591, 25'd2760}, '{25'd1971, 25'd5322, 25'd1380, 25'd5322, 25'd1183}, '{25'd5914, 25'd4731, 25'd1774, 25'd1971, 25'd4731}, '{25'd5125, 25'd3548, 25'd2168, 25'd1577, 25'd1183}}, '{'{25'd5717, 25'd6505, 25'd2168, 25'd3548, 25'd4731}, '{25'd3745, 25'd3351, 25'd3943, 25'd1774, 25'd789}, '{25'd7097, 25'd7491, 25'd3943, 25'd3351, 25'd4731}, '{25'd4731, 25'd5914, 25'd2957, 25'd4534, 25'd3154}, '{25'd8477, 25'd4928, 25'd7097, 25'd4928, 25'd3351}}, '{'{25'd6900, 25'd19319, 25'd25035, 25'd14982, 25'd13405}, '{25'd591, 25'd10054, 25'd19516, 25'd8082, 25'd12616}, '{25'd19910, 25'd23458, 25'd25035, 25'd24641, 25'd25035}, '{25'd9856, 25'd18136, 25'd21093, 25'd12813, 25'd13996}, '{-25'd3351, 25'd7885, 25'd8477, 25'd4140, 25'd2366}}, '{'{25'd1380, 25'd1971, -25'd197, -25'd986, 25'd2957}, '{-25'd1183, 25'd2563, -25'd197, 25'd2760, 25'd986}, '{25'd2957, 25'd2366, 25'd0, -25'd1183, -25'd986}, '{25'd1971, -25'd789, -25'd986, 25'd2760, 25'd1577}, '{-25'd789, 25'd2563, 25'd986, -25'd197, -25'd1577}}, '{'{-25'd4928, -25'd2366, -25'd394, -25'd3943, -25'd5322}, '{-25'd2366, -25'd4731, -25'd3548, -25'd1183, -25'd4731}, '{-25'd1774, -25'd789, -25'd986, -25'd4731, -25'd1971}, '{-25'd1380, -25'd2168, -25'd4928, -25'd4337, -25'd2563}, '{-25'd986, -25'd3154, -25'd1183, -25'd1380, -25'd3745}}, '{'{25'd1971, 25'd2366, 25'd2563, 25'd3154, 25'd2168}, '{25'd1774, 25'd789, -25'd986, 25'd2168, -25'd197}, '{-25'd591, 25'd2957, 25'd986, -25'd591, -25'd1380}, '{25'd2168, 25'd2760, 25'd1577, 25'd986, -25'd986}, '{25'd1774, -25'd1380, -25'd1380, -25'd591, 25'd591}}, '{'{25'd12025, 25'd9462, 25'd14588, 25'd14193, 25'd14588}, '{25'd14193, 25'd12419, 25'd11828, 25'd13208, 25'd11236}, '{25'd11828, 25'd12813, 25'd11828, 25'd9856, 25'd10251}, '{25'd10448, 25'd12025, 25'd11236, 25'd13996, 25'd11631}, '{25'd10645, 25'd11433, 25'd12813, 25'd12616, 25'd11828}}, '{'{25'd4731, 25'd2168, 25'd5717, 25'd1183, 25'd5322}, '{25'd5322, 25'd3943, 25'd3943, 25'd4731, 25'd4534}, '{25'd1971, 25'd2366, 25'd789, 25'd2957, 25'd1577}, '{25'd2563, 25'd2760, 25'd5322, 25'd1183, 25'd3943}, '{25'd1774, 25'd3548, 25'd3351, 25'd1380, 25'd5717}}, '{'{-25'd197, 25'd591, 25'd3943, 25'd1774, 25'd591}, '{-25'd394, 25'd3745, 25'd2957, 25'd1183, 25'd986}, '{25'd394, 25'd1971, 25'd2760, 25'd2168, 25'd197}, '{25'd197, 25'd3154, 25'd2563, 25'd2168, 25'd789}, '{25'd2366, 25'd1380, -25'd394, 25'd591, 25'd2957}}, '{'{25'd2957, 25'd4534, 25'd3548, 25'd2760, 25'd3943}, '{25'd6308, 25'd6308, 25'd1577, 25'd1183, 25'd4731}, '{25'd5125, 25'd2168, 25'd3745, 25'd4534, 25'd5520}, '{25'd2168, 25'd1971, 25'd4337, 25'd2366, 25'd6702}, '{25'd1380, 25'd3548, 25'd4928, 25'd2957, 25'd6111}}, '{'{25'd1971, 25'd1183, 25'd986, 25'd1577, 25'd1577}, '{25'd986, 25'd0, -25'd591, 25'd0, 25'd2563}, '{25'd1380, 25'd1577, 25'd3154, 25'd1183, -25'd394}, '{25'd2563, 25'd197, 25'd2957, -25'd197, 25'd2168}, '{25'd2563, -25'd1380, 25'd2760, 25'd1380, 25'd2366}}, '{'{25'd2168, -25'd986, -25'd591, 25'd2563, 25'd197}, '{-25'd789, -25'd1183, 25'd197, 25'd789, -25'd986}, '{25'd1971, 25'd3351, 25'd3154, 25'd2957, 25'd1774}, '{25'd1183, 25'd2366, 25'd197, -25'd1380, 25'd0}, '{-25'd1183, 25'd1183, -25'd394, 25'd394, 25'd3548}}, '{'{25'd6702, 25'd5322, 25'd4928, 25'd5914, 25'd1774}, '{25'd5717, 25'd2760, 25'd986, 25'd2366, 25'd3351}, '{25'd6111, 25'd5914, 25'd2760, 25'd2563, 25'd1774}, '{25'd5520, 25'd2957, 25'd1971, 25'd789, 25'd5125}, '{25'd2563, 25'd1183, 25'd4140, 25'd5322, 25'd6505}}, '{'{25'd4534, 25'd1380, 25'd6505, 25'd5520, 25'd3943}, '{25'd3154, 25'd5717, 25'd6900, 25'd3745, 25'd5520}, '{25'd6308, 25'd3548, 25'd4337, 25'd5520, 25'd8477}, '{25'd5322, 25'd3745, 25'd6505, 25'd6900, 25'd7097}, '{25'd5717, 25'd3548, 25'd5914, 25'd6900, 25'd9068}}, '{'{25'd2563, 25'd789, 25'd1183, 25'd3745, 25'd7491}, '{25'd3154, 25'd1971, 25'd5125, 25'd5717, 25'd8279}, '{25'd3943, 25'd5717, 25'd2760, 25'd3943, 25'd6308}, '{25'd3351, 25'd2760, 25'd5125, 25'd2957, 25'd6505}, '{25'd5717, 25'd4140, 25'd3154, 25'd1380, 25'd4731}}, '{'{-25'd3745, -25'd4534, -25'd1183, -25'd2957, -25'd394}, '{-25'd2760, -25'd3745, -25'd2563, 25'd0, -25'd3548}, '{-25'd789, -25'd3154, -25'd3154, -25'd4337, -25'd4534}, '{-25'd591, -25'd1774, -25'd2168, -25'd4731, -25'd3154}, '{-25'd4731, -25'd2366, -25'd2760, -25'd4731, -25'd2168}}, '{'{25'd24444, 25'd23655, 25'd20699, 25'd20107, 25'd16953}, '{25'd19122, 25'd19319, 25'd20896, 25'd18333, 25'd14982}, '{25'd17742, 25'd18727, 25'd19122, 25'd15770, 25'd12813}, '{25'd15573, 25'd15967, 25'd17150, 25'd12813, 25'd11236}, '{25'd19319, 25'd18530, 25'd19516, 25'd17347, 25'd14588}}, '{'{25'd13011, 25'd12616, 25'd13799, 25'd10842, 25'd10645}, '{25'd12813, 25'd12222, 25'd10251, 25'd9265, 25'd9659}, '{25'd15967, 25'd13208, 25'd13405, 25'd10054, 25'd10054}, '{25'd12813, 25'd11039, 25'd11828, 25'd10645, 25'd9856}, '{25'd13799, 25'd10842, 25'd11433, 25'd11631, 25'd14193}}, '{'{25'd3745, 25'd986, 25'd3548, 25'd2957, 25'd3351}, '{25'd1183, 25'd3943, 25'd2563, 25'd1577, 25'd3745}, '{25'd2563, 25'd2168, -25'd197, 25'd3745, 25'd2168}, '{25'd986, -25'd197, -25'd197, 25'd5125, 25'd3548}, '{25'd4928, 25'd1971, 25'd2168, 25'd6505, 25'd5520}}, '{'{-25'd4140, 25'd394, 25'd394, -25'd197, 25'd1380}, '{25'd15770, 25'd18136, 25'd18727, 25'd16953, 25'd19319}, '{25'd16953, 25'd20896, 25'd19910, 25'd18924, 25'd24444}, '{25'd11631, 25'd10448, 25'd18136, 25'd17150, 25'd20304}, '{25'd8871, 25'd7097, 25'd10842, 25'd12813, 25'd15376}}, '{'{25'd13996, 25'd13208, 25'd9462, 25'd10842, 25'd10251}, '{25'd10054, 25'd11236, 25'd12222, 25'd8082, 25'd8674}, '{25'd8477, 25'd10251, 25'd7688, 25'd10251, 25'd11433}, '{25'd8082, 25'd6505, 25'd9856, 25'd8871, 25'd9856}, '{25'd11828, 25'd11039, 25'd7688, 25'd8871, 25'd10054}}, '{'{25'd6702, 25'd6505, 25'd5717, 25'd5520, 25'd7688}, '{25'd7688, 25'd4928, 25'd5717, 25'd9462, 25'd8279}, '{25'd8674, 25'd6702, 25'd8871, 25'd9856, 25'd7294}, '{25'd9659, 25'd8477, 25'd5717, 25'd6505, 25'd12419}, '{25'd12222, 25'd11631, 25'd10842, 25'd12616, 25'd11828}}, '{'{25'd11236, 25'd10054, 25'd10054, 25'd13011, 25'd11828}, '{25'd10448, 25'd10251, 25'd11433, 25'd10251, 25'd11433}, '{25'd10251, 25'd8477, 25'd8674, 25'd9265, 25'd11828}, '{25'd14588, 25'd10842, 25'd12616, 25'd11433, 25'd10645}, '{25'd12813, 25'd13011, 25'd14390, 25'd13602, 25'd10448}}, '{'{25'd12813, 25'd9265, 25'd11828, 25'd10054, 25'd11828}, '{25'd10251, 25'd12025, 25'd9462, 25'd7294, 25'd9856}, '{25'd9068, 25'd8477, 25'd11236, 25'd10842, 25'd8871}, '{25'd10251, 25'd11433, 25'd7294, 25'd10251, 25'd8871}, '{25'd10842, 25'd11236, 25'd11236, 25'd7491, 25'd9659}}, '{'{25'd2366, 25'd3548, 25'd2957, 25'd789, 25'd3351}, '{25'd1774, 25'd2760, 25'd3154, 25'd394, 25'd789}, '{25'd3943, 25'd1183, 25'd1774, -25'd394, 25'd3548}, '{25'd2563, -25'd197, 25'd197, 25'd394, 25'd4928}, '{25'd591, -25'd197, 25'd2366, 25'd1971, 25'd3351}}, '{'{25'd3943, 25'd2168, 25'd4928, 25'd4140, 25'd4731}, '{25'd1183, 25'd3351, 25'd5322, 25'd6505, 25'd6900}, '{25'd5914, 25'd1380, 25'd5322, 25'd6702, 25'd7491}, '{25'd6505, 25'd5520, 25'd5322, 25'd7294, 25'd7688}, '{25'd6111, 25'd5125, 25'd5717, 25'd3548, 25'd4534}}, '{'{25'd2957, 25'd2760, 25'd394, 25'd2760, 25'd2957}, '{25'd789, -25'd197, 25'd1774, -25'd591, 25'd2168}, '{-25'd394, -25'd986, -25'd591, 25'd3548, 25'd2168}, '{25'd1774, 25'd2366, 25'd197, 25'd2957, 25'd2957}, '{25'd1380, 25'd2760, 25'd2957, -25'd197, -25'd197}}, '{'{25'd8674, 25'd4731, 25'd3351, 25'd2563, 25'd7294}, '{25'd8871, 25'd3154, 25'd2168, 25'd5520, 25'd3745}, '{25'd5322, 25'd3943, 25'd3943, 25'd3351, 25'd5125}, '{25'd3943, 25'd6505, 25'd6308, 25'd6111, 25'd2957}, '{25'd5125, 25'd3548, 25'd2563, 25'd2760, 25'd3943}}, '{'{25'd12222, 25'd11039, 25'd10645, 25'd17939, 25'd16559}, '{25'd12813, 25'd7294, 25'd12419, 25'd16953, 25'd16165}, '{25'd7491, 25'd6702, 25'd10842, 25'd13996, 25'd16756}, '{25'd10842, 25'd8674, 25'd13405, 25'd13799, 25'd18530}, '{25'd12419, 25'd11236, 25'd16756, 25'd18333, 25'd18333}}},
    '{'{'{-25'd1191, -25'd198, 25'd2382, 25'd3572, -25'd198}, '{25'd794, 25'd2382, -25'd794, 25'd794, 25'd1191}, '{25'd3771, 25'd2779, 25'd2977, 25'd2779, -25'd595}, '{25'd794, 25'd1588, -25'd595, 25'd3969, 25'd1191}, '{25'd3175, 25'd0, 25'd3572, -25'd794, 25'd3374}}, '{'{25'd6946, 25'd6351, 25'd3572, 25'd2977, 25'd6549}, '{25'd4565, 25'd6946, 25'd6351, 25'd1786, 25'd2779}, '{25'd3771, 25'd4168, 25'd4565, 25'd2580, 25'd4565}, '{25'd6152, 25'd3175, 25'd1588, 25'd5557, 25'd3572}, '{25'd4168, 25'd4366, 25'd3175, 25'd7939, 25'd5359}}, '{'{25'd1985, -25'd397, 25'd2580, 25'd2977, 25'd1389}, '{25'd2977, 25'd2779, 25'd198, 25'd1786, -25'd1191}, '{25'd2977, 25'd198, 25'd992, 25'd3175, 25'd595}, '{-25'd595, -25'd198, 25'd3374, 25'd1588, -25'd198}, '{-25'd198, 25'd198, 25'd2183, 25'd2977, 25'd1389}}, '{'{25'd2183, 25'd3374, 25'd4168, 25'd4366, 25'd2580}, '{25'd3572, 25'd2779, 25'd2382, 25'd3771, 25'd2779}, '{25'd1786, 25'd3771, 25'd3771, 25'd2779, 25'd3969}, '{25'd3969, 25'd2779, 25'd5557, 25'd1191, 25'd2580}, '{25'd5557, 25'd1389, 25'd2779, 25'd1389, 25'd595}}, '{'{25'd5756, 25'd5954, 25'd3969, 25'd1786, 25'd4168}, '{25'd4962, 25'd2183, 25'd2977, 25'd2779, 25'd3374}, '{25'd6152, 25'd6152, 25'd6152, 25'd4168, 25'd1985}, '{25'd4962, 25'd5954, 25'd2977, 25'd2183, 25'd5756}, '{25'd8931, 25'd7343, 25'd3771, 25'd3771, 25'd6748}}, '{'{25'd2977, 25'd21236, 25'd25205, 25'd13297, 25'd13099}, '{-25'd3771, 25'd10717, 25'd20442, 25'd7343, 25'd7343}, '{25'd11114, 25'd16671, 25'd21236, 25'd14091, 25'd17267}, '{25'd10717, 25'd17267, 25'd22228, 25'd13694, 25'd14488}, '{25'd1985, 25'd10320, 25'd14686, 25'd992, 25'd6351}}, '{'{25'd2382, 25'd2580, 25'd2382, -25'd1588, -25'd992}, '{25'd1786, -25'd2183, -25'd1588, -25'd397, 25'd3175}, '{25'd2382, 25'd0, -25'd1985, 25'd1985, 25'd2779}, '{-25'd992, 25'd1786, 25'd1389, -25'd794, -25'd595}, '{25'd595, 25'd1389, 25'd992, -25'd794, 25'd198}}, '{'{-25'd3771, -25'd2382, -25'd794, -25'd3771, -25'd1588}, '{-25'd3374, -25'd3969, -25'd1985, -25'd198, -25'd1985}, '{-25'd992, -25'd2580, -25'd3572, -25'd2580, -25'd595}, '{-25'd1588, -25'd1985, -25'd2382, -25'd4962, -25'd4565}, '{-25'd4962, -25'd3175, -25'd397, -25'd4565, -25'd3175}}, '{'{-25'd1191, 25'd2580, 25'd2779, 25'd595, 25'd2580}, '{25'd1389, 25'd2382, 25'd1985, -25'd595, 25'd2183}, '{25'd2580, 25'd2183, -25'd794, 25'd1588, -25'd595}, '{-25'd992, 25'd1389, 25'd2183, -25'd1191, 25'd1191}, '{25'd1191, 25'd2580, 25'd2977, -25'd1588, -25'd794}}, '{'{25'd12702, 25'd12900, 25'd10916, 25'd11908, 25'd10916}, '{25'd16274, 25'd11511, 25'd9923, 25'd11908, 25'd14091}, '{25'd13297, 25'd10122, 25'd11709, 25'd14686, 25'd11114}, '{25'd13893, 25'd10519, 25'd11511, 25'd14091, 25'd13893}, '{25'd13694, 25'd8336, 25'd13893, 25'd9526, 25'd10916}}, '{'{25'd794, 25'd1588, 25'd4962, 25'd4366, 25'd1588}, '{25'd3771, 25'd1191, 25'd4763, 25'd2779, 25'd4763}, '{25'd2779, 25'd3771, 25'd4962, 25'd4168, 25'd4565}, '{25'd3771, 25'd992, 25'd4763, 25'd2580, 25'd1389}, '{25'd2779, 25'd3969, 25'd992, 25'd2382, 25'd5557}}, '{'{-25'd595, 25'd794, 25'd1191, 25'd198, 25'd1191}, '{25'd2382, 25'd992, 25'd3771, 25'd397, 25'd3374}, '{25'd1588, 25'd2183, 25'd2977, 25'd4168, 25'd1786}, '{25'd2183, 25'd2580, -25'd198, 25'd3572, 25'd1786}, '{25'd2779, 25'd1389, 25'd2977, 25'd397, 25'd1191}}, '{'{25'd6351, 25'd4366, 25'd4763, 25'd1985, 25'd3175}, '{25'd1389, 25'd1985, 25'd5359, 25'd4366, 25'd3175}, '{25'd4962, 25'd2382, 25'd4366, 25'd1588, 25'd3572}, '{25'd2382, 25'd1786, 25'd5359, 25'd2382, 25'd5954}, '{25'd5557, 25'd5359, 25'd1985, 25'd7343, 25'd5160}}, '{'{-25'd595, 25'd1588, -25'd794, 25'd1786, -25'd992}, '{25'd1588, 25'd0, 25'd1588, 25'd1588, 25'd397}, '{-25'd397, 25'd198, -25'd397, 25'd2382, 25'd3175}, '{-25'd794, 25'd198, 25'd397, 25'd2977, 25'd1786}, '{25'd198, 25'd1389, -25'd397, 25'd3374, -25'd794}}, '{'{25'd1389, 25'd595, 25'd1588, 25'd2382, 25'd2580}, '{25'd1588, 25'd2580, 25'd1786, 25'd1588, 25'd1588}, '{25'd595, 25'd2183, 25'd992, 25'd2183, -25'd198}, '{-25'd397, 25'd198, -25'd1191, 25'd2580, 25'd2580}, '{25'd3175, -25'd1588, 25'd0, 25'd198, 25'd992}}, '{'{25'd7542, 25'd3572, 25'd2779, 25'd2580, 25'd4565}, '{25'd7740, 25'd4366, 25'd3175, 25'd397, 25'd992}, '{25'd6748, 25'd3572, 25'd3771, 25'd3771, 25'd3374}, '{25'd6152, 25'd3771, 25'd397, 25'd2779, 25'd4565}, '{25'd2977, 25'd4763, 25'd2382, 25'd4565, 25'd7145}}, '{'{25'd1985, 25'd3572, 25'd2779, 25'd3175, 25'd3175}, '{25'd4366, 25'd5160, 25'd7542, 25'd5954, 25'd4168}, '{25'd8336, 25'd6748, 25'd4366, 25'd7542, 25'd5557}, '{25'd6152, 25'd5756, 25'd8534, 25'd5954, 25'd4763}, '{25'd5954, 25'd5756, 25'd4962, 25'd4962, 25'd6152}}, '{'{25'd794, 25'd2779, 25'd5756, 25'd6351, 25'd6152}, '{25'd2977, 25'd2183, 25'd4962, 25'd3771, 25'd7740}, '{25'd2977, 25'd4168, 25'd2779, 25'd5557, 25'd2779}, '{25'd2779, 25'd2779, 25'd3572, 25'd1786, 25'd6152}, '{25'd4565, 25'd5359, 25'd3771, 25'd1191, 25'd1786}}, '{'{-25'd2183, -25'd2779, -25'd4565, -25'd595, -25'd1985}, '{-25'd3572, -25'd3175, -25'd3175, 25'd0, -25'd2977}, '{-25'd198, -25'd4565, -25'd3771, -25'd3969, -25'd1985}, '{-25'd3969, -25'd2779, -25'd4565, -25'd992, -25'd4763}, '{-25'd198, -25'd992, -25'd3771, -25'd2977, -25'd4366}}, '{'{25'd23022, 25'd25007, 25'd20640, 25'd18259, 25'd14488}, '{25'd24808, 25'd22228, 25'd17663, 25'd16076, 25'd14686}, '{25'd20243, 25'd19648, 25'd17267, 25'd14290, 25'd8732}, '{25'd19251, 25'd15083, 25'd18457, 25'd14290, 25'd11908}, '{25'd18457, 25'd17862, 25'd16473, 25'd17068, 25'd11114}}, '{'{25'd14488, 25'd13694, 25'd11313, 25'd10122, 25'd10122}, '{25'd13297, 25'd9129, 25'd12702, 25'd9129, 25'd13297}, '{25'd11114, 25'd11511, 25'd12702, 25'd8931, 25'd9328}, '{25'd10717, 25'd12503, 25'd10916, 25'd10519, 25'd14091}, '{25'd12106, 25'd10122, 25'd11313, 25'd10519, 25'd13496}}, '{'{25'd3771, 25'd2382, 25'd1191, 25'd4962, 25'd2580}, '{25'd1985, 25'd2580, 25'd1191, -25'd397, 25'd992}, '{-25'd595, 25'd1389, 25'd2183, 25'd2183, 25'd1588}, '{25'd3175, 25'd3374, 25'd1389, 25'd992, 25'd4962}, '{25'd3771, 25'd4565, 25'd4962, 25'd5954, 25'd4962}}, '{'{-25'd2977, -25'd1588, 25'd7740, -25'd198, 25'd1588}, '{25'd11114, 25'd13893, 25'd17465, 25'd12702, 25'd16870}, '{25'd16076, 25'd19847, 25'd22030, 25'd20640, 25'd24411}, '{25'd9129, 25'd11511, 25'd19648, 25'd19053, 25'd21037}, '{25'd5359, 25'd5954, 25'd15282, 25'd12106, 25'd19053}}, '{'{25'd12900, 25'd9328, 25'd12503, 25'd12305, 25'd8336}, '{25'd10519, 25'd12900, 25'd11511, 25'd11114, 25'd9923}, '{25'd10320, 25'd9725, 25'd7740, 25'd8931, 25'd11709}, '{25'd7939, 25'd10916, 25'd7343, 25'd6748, 25'd11114}, '{25'd9923, 25'd9923, 25'd10717, 25'd8931, 25'd6748}}, '{'{25'd6351, 25'd5359, 25'd6351, 25'd7145, 25'd5160}, '{25'd6748, 25'd4763, 25'd6946, 25'd4366, 25'd5160}, '{25'd8336, 25'd7740, 25'd9129, 25'd10320, 25'd8534}, '{25'd12106, 25'd7939, 25'd8732, 25'd12305, 25'd9328}, '{25'd11908, 25'd10916, 25'd13099, 25'd10916, 25'd10717}}, '{'{25'd10122, 25'd11908, 25'd8732, 25'd12702, 25'd10916}, '{25'd12503, 25'd10320, 25'd11114, 25'd8732, 25'd10122}, '{25'd12702, 25'd8137, 25'd11511, 25'd12305, 25'd11908}, '{25'd13694, 25'd10916, 25'd12106, 25'd11114, 25'd10320}, '{25'd14488, 25'd11313, 25'd12503, 25'd10916, 25'd11114}}, '{'{25'd11709, 25'd10122, 25'd12305, 25'd9725, 25'd8137}, '{25'd12305, 25'd8137, 25'd10916, 25'd8931, 25'd10916}, '{25'd11114, 25'd8534, 25'd8137, 25'd10717, 25'd9328}, '{25'd11908, 25'd9526, 25'd7740, 25'd7939, 25'd10916}, '{25'd12106, 25'd10320, 25'd9526, 25'd10122, 25'd8732}}, '{'{25'd3771, -25'd198, 25'd397, 25'd397, 25'd1588}, '{25'd2779, 25'd3771, -25'd397, 25'd1389, 25'd4168}, '{25'd2977, 25'd3374, 25'd992, 25'd2382, 25'd2779}, '{25'd1191, -25'd198, 25'd992, 25'd1389, 25'd3374}, '{25'd2779, 25'd2779, 25'd3771, 25'd3771, 25'd5359}}, '{'{25'd5160, 25'd4168, 25'd2580, 25'd3771, 25'd5359}, '{25'd1786, 25'd4763, 25'd4763, 25'd7145, 25'd7939}, '{25'd5954, 25'd3374, 25'd3771, 25'd5954, 25'd3771}, '{25'd3771, 25'd4565, 25'd5160, 25'd3969, 25'd5160}, '{25'd6748, 25'd4565, 25'd3969, 25'd7939, 25'd8336}}, '{'{25'd992, -25'd1389, 25'd2183, 25'd3175, 25'd3374}, '{25'd2977, -25'd595, -25'd992, 25'd2183, 25'd3572}, '{25'd2779, 25'd992, -25'd198, 25'd198, 25'd3374}, '{25'd2382, 25'd3175, 25'd2779, -25'd397, -25'd397}, '{25'd3175, 25'd1191, 25'd1786, -25'd595, 25'd3771}}, '{'{25'd8137, 25'd4366, 25'd5160, 25'd3374, 25'd4168}, '{25'd7145, 25'd3969, 25'd3572, 25'd5160, 25'd4763}, '{25'd4763, 25'd5756, 25'd2183, 25'd2779, 25'd4168}, '{25'd3969, 25'd6549, 25'd3771, 25'd5557, 25'd4168}, '{25'd4763, 25'd3175, 25'd6946, 25'd3374, 25'd3572}}, '{'{25'd12106, 25'd10916, 25'd12702, 25'd17068, 25'd20243}, '{25'd9526, 25'd6946, 25'd10122, 25'd16076, 25'd18457}, '{25'd9923, 25'd9328, 25'd12900, 25'd15679, 25'd14686}, '{25'd9328, 25'd8732, 25'd13893, 25'd13297, 25'd15083}, '{25'd14091, 25'd13297, 25'd14091, 25'd15877, 25'd17068}}}
};
