localparam bit signed [0:2][35:0] Bias3 = '{36'd0, 36'd0, 36'd0};
