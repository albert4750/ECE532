localparam bit signed [0:63][47:0] Bias1 = '{48'd2656677, 48'd1113730, 48'd3027799, -48'd2889267, -48'd2267660, 48'd1350262, -48'd2729511, -48'd3393636, 48'd433726, -48'd4461216, -48'd783634, 48'd2073061, 48'd3691289, -48'd535444, 48'd2023121, -48'd777857, -48'd466149, -48'd3266590, 48'd264985, 48'd1073415, 48'd764155, 48'd1437437, 48'd3575592, -48'd3203198, -48'd3867110, 48'd909309, -48'd630225, -48'd1892020, -48'd2500874, 48'd2073900, 48'd2958129, -48'd392867, 48'd2621255, -48'd1566216, 48'd251271, -48'd556158, 48'd3538772, -48'd2039337, 48'd4246514, 48'd1850222, -48'd1960709, -48'd1193555, 48'd1450934, -48'd3840564, 48'd2391534, 48'd2063727, -48'd2082220, -48'd1934319, -48'd7612231, 48'd757458, -48'd4264268, -48'd2324221, -48'd498146, 48'd3496729, 48'd220376, -48'd208004, 48'd130498, -48'd2744673, 48'd4319400, -48'd6067323, 48'd3499428, 48'd1480624, 48'd6083084, 48'd739223};
