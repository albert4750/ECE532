localparam bit signed [0:7][0:7][0:2][0:2][19:0] Weight2 = '{
    '{'{'{-20'd91392, -20'd67200, -20'd72576}, '{-20'd131713, -20'd118273, -20'd231169}, '{20'd107520, -20'd5376, -20'd80640}}, '{'{20'd2688, -20'd24192, 20'd24192}, '{20'd32256, -20'd5376, 20'd18816}, '{20'd21504, 20'd21504, 20'd45696}}, '{'{20'd129025, 20'd102144, -20'd215041}, '{20'd142465, 20'd118273, 20'd145153}, '{-20'd147841, 20'd161281, 20'd301057}}, '{'{-20'd174721, 20'd59136, -20'd29568}, '{20'd10752, 20'd341378, 20'd180097}, '{-20'd110208, 20'd45696, -20'd142465}}, '{'{20'd61824, 20'd53760, 20'd67200}, '{20'd8064, 20'd10752, 20'd64512}, '{20'd75264, 20'd34944, 20'd26880}}, '{'{20'd53760, 20'd43008, 20'd18816}, '{-20'd180097, -20'd8064, -20'd158593}, '{20'd5376, 20'd120961, -20'd37632}}, '{'{-20'd94080, 20'd180097, 20'd24192}, '{-20'd2688, 20'd147841, 20'd94080}, '{-20'd18816, 20'd110208, -20'd2688}}, '{'{-20'd96768, 20'd88704, 20'd53760}, '{-20'd56448, -20'd40320, 20'd104832}, '{-20'd2688, 20'd43008, 20'd8064}}},
    '{'{'{-20'd118974, -20'd114800, -20'd25047}, '{-20'd128367, -20'd76185, -20'd83491}, '{-20'd76185, -20'd61574, -20'd13567}}, '{'{20'd0, -20'd27135, 20'd77229}, '{20'd13567, -20'd38614, -20'd43833}, '{-20'd67836, 20'd59487, 20'd30265}}, '{'{-20'd19829, -20'd2087, -20'd10436}, '{-20'd5218, 20'd29222, -20'd75142}, '{20'd132542, -20'd74098, -20'd77229}}, '{'{-20'd97058, 20'd0, -20'd70967}, '{-20'd90796, -20'd27135, 20'd2087}, '{-20'd81404, 20'd75142, -20'd89753}}, '{'{-20'd29222, -20'd75142, -20'd49051}, '{20'd41745, 20'd19829, 20'd40702}, '{-20'd58444, 20'd21916, 20'd81404}}, '{'{20'd38614, -20'd61574, -20'd74098}, '{20'd98102, -20'd65749, -20'd76185}, '{20'd29222, -20'd64705, 20'd28178}}, '{'{-20'd20873, -20'd112713, -20'd45920}, '{-20'd32353, 20'd0, -20'd75142}, '{-20'd102276, -20'd110625, -20'd68880}}, '{'{20'd11480, -20'd57400, -20'd101233}, '{-20'd11480, -20'd81404, 20'd8349}, '{-20'd9393, -20'd50094, -20'd55313}}},
    '{'{'{20'd2301, -20'd214015, -20'd64435}, '{-20'd253136, -20'd101255, 20'd174894}, '{20'd48326, 20'd73640, 20'd200208}}, '{'{20'd34519, 20'd128869, 20'd46025}, '{20'd131171, 20'd46025, -20'd29916}, '{20'd124267, 20'd64435, 20'd96652}}, '{'{-20'd82845, -20'd69037, -20'd52929}, '{-20'd32217, 20'd124267, 20'd57531}, '{-20'd18410, 20'd101255, 20'd62133}}, '{'{-20'd269245, 20'd151882, -20'd6904}, '{20'd227823, 20'd292258, 20'd292258}, '{-20'd191003, 20'd126568, -20'd105857}}, '{'{20'd64435, 20'd29916, 20'd9205}, '{20'd115062, 20'd119665, 20'd108158}, '{20'd92050, -20'd13807, 20'd69037}}, '{'{20'd98953, 20'd23012, 20'd131171}, '{-20'd105857, -20'd294559, -20'd135773}, '{20'd23012, 20'd4602, -20'd50627}}, '{'{20'd13807, 20'd156484, 20'd140376}, '{20'd25314, 20'd117363, -20'd11506}, '{20'd62133, 20'd2301, 20'd80543}}, '{'{20'd52929, -20'd9205, 20'd50627}, '{20'd112761, 20'd165689, 20'd89748}, '{-20'd98953, -20'd41422, -20'd29916}}},
    '{'{'{-20'd52772, -20'd50259, 20'd158317}, '{-20'd268887, -20'd140726, 20'd238732}, '{-20'd160830, -20'd115596, -20'd243758}}, '{'{-20'd42720, 20'd32669, 20'd95493}, '{20'd7539, 20'd98006, 20'd123135}, '{20'd35182, 20'd113083, -20'd40207}}, '{'{-20'd85441, 20'd82928, -20'd135700}, '{-20'd2513, 20'd25130, -20'd55285}, '{-20'd35182, 20'd87954, 20'd319147}}, '{'{-20'd55285, 20'd211089, 20'd87954}, '{-20'd77902, 20'd196011, 20'd173395}, '{-20'd233706, -20'd50259, 20'd2513}}, '{'{20'd105545, 20'd92980, 20'd42720}, '{20'd12565, 20'd37694, 20'd67850}, '{20'd115596, 20'd27643, 20'd12565}}, '{'{20'd128161, -20'd236219, 20'd17591}, '{-20'd118109, -20'd180933, -20'd17591}, '{-20'd40207, -20'd42720, -20'd130674}}, '{'{20'd20104, -20'd42720, -20'd62824}, '{20'd135700, -20'd45233, 20'd37694}, '{-20'd17591, 20'd110570, 20'd57798}}, '{'{20'd85441, 20'd82928, 20'd185959}, '{20'd241245, 20'd72876, 20'd15078}, '{20'd17591, 20'd20104, 20'd55285}}},
    '{'{'{-20'd102483, -20'd31607, -20'd67045}, '{-20'd5747, -20'd120681, -20'd3831}, '{-20'd122596, -20'd28734, -20'd13409}}, '{'{-20'd13409, -20'd2873, -20'd52678}, '{-20'd14367, -20'd68960, 20'd958}, '{-20'd102483, 20'd17240, -20'd12451}}, '{'{-20'd38311, -20'd109187, -20'd97694}, '{-20'd35438, -20'd38311, 20'd34480}, '{-20'd24902, 20'd40227, 20'd38311}}, '{'{-20'd12451, -20'd20113, -20'd19156}, '{20'd10536, -20'd118765, -20'd22987}, '{-20'd75665, -20'd6704, -20'd42143}}, '{'{-20'd52678, -20'd77581, -20'd9578}, '{20'd28734, -20'd55552, -20'd100567}, '{-20'd28734, 20'd20113, -20'd16282}}, '{'{-20'd1916, -20'd93863, -20'd80454}, '{20'd13409, -20'd51720, -20'd25860}, '{-20'd45016, 20'd3831, 20'd22987}}, '{'{-20'd68960, -20'd87158, -20'd119723}, '{-20'd33522, 20'd19156, -20'd55552}, '{-20'd48847, 20'd10536, -20'd75665}}, '{'{20'd28734, -20'd56509, 20'd19156}, '{-20'd113976, -20'd51720, -20'd108230}, '{-20'd101525, -20'd39269, -20'd73749}}},
    '{'{'{-20'd125861, 20'd32364, -20'd38358}, '{-20'd153430, -20'd116271, 20'd29967}, '{-20'd20377, 20'd4795, 20'd69523}}, '{'{-20'd19179, 20'd11987, 20'd34762}, '{-20'd15583, -20'd76715, -20'd11987}, '{20'd14384, -20'd14384, 20'd9589}}, '{'{20'd29967, 20'd39556, 20'd45550}, '{-20'd11987, 20'd53940, 20'd55139}, '{-20'd2397, -20'd5993, -20'd39556}}, '{'{-20'd5993, 20'd46748, -20'd57536}, '{-20'd131854, 20'd74318, -20'd58735}, '{20'd22775, 20'd97093, -20'd52742}}, '{'{-20'd83907, -20'd59934, 20'd8391}, '{-20'd21576, -20'd28768, -20'd99490}, '{-20'd117470, -20'd116271, -20'd49146}}, '{'{-20'd41954, -20'd38358, 20'd11987}, '{-20'd89900, -20'd73119, -20'd82708}, '{-20'd15583, -20'd7192, -20'd106682}}, '{'{-20'd43152, 20'd0, -20'd89900}, '{-20'd59934, -20'd80311, -20'd64728}, '{-20'd94695, -20'd107881, -20'd47947}}, '{'{20'd31166, -20'd4795, -20'd98291}, '{20'd52742, -20'd93497, -20'd13185}, '{20'd53940, -20'd45550, -20'd29967}}},
    '{'{'{20'd13344, 20'd48291, 20'd59093}, '{-20'd8896, -20'd50197, 20'd33676}, '{-20'd17156, -20'd61634, 20'd55280}}, '{'{-20'd3812, 20'd51468, -20'd47655}, '{-20'd43843, 20'd635, 20'd2542}, '{20'd52103, -20'd49562, 20'd635}}, '{'{-20'd81332, 20'd69895, 20'd2542}, '{20'd26687, 20'd60363, -20'd20333}, '{20'd63541, -20'd11437, 20'd73072}}, '{'{20'd57822, -20'd76249, -20'd44478}, '{20'd6989, -20'd75613, 20'd6989}, '{-20'd72436, 20'd19698, -20'd34312}}, '{'{-20'd41301, -20'd17791, -20'd63541}, '{20'd54009, -20'd57186, -20'd27322}, '{-20'd17791, -20'd46385, 20'd45114}}, '{'{-20'd70530, -20'd28593, 20'd12708}, '{-20'd22875, 20'd17156, -20'd22875}, '{20'd15885, -20'd12708, -20'd64811}}, '{'{-20'd31135, -20'd79426, -20'd38760}, '{-20'd72436, -20'd4448, -20'd61634}, '{-20'd15250, -20'd72436, -20'd74978}}, '{'{-20'd57822, -20'd1906, -20'd635}, '{20'd60363, -20'd65447, -20'd38760}, '{20'd59728, -20'd78790, -20'd65447}}},
    '{'{'{-20'd46438, -20'd78016, -20'd36221}, '{-20'd31578, 20'd19504, -20'd27863}, '{-20'd76158, -20'd46438, -20'd52010}}, '{'{-20'd84517, -20'd104949, 20'd32506}, '{20'd0, 20'd23219, -20'd115166}, '{-20'd48295, -20'd34364, 20'd24148}}, '{'{20'd14860, -20'd74300, -20'd76158}, '{-20'd117023, -20'd70585, 20'd29720}, '{-20'd10216, 20'd36221, 20'd13003}}, '{'{-20'd37150, -20'd6501, -20'd19504}, '{-20'd104021, 20'd39008, 20'd33435}, '{-20'd48295, 20'd39937, -20'd48295}}, '{'{20'd39937, 20'd25076, -20'd16718}, '{-20'd48295, 20'd31578, -20'd64084}, '{20'd35293, 20'd8359, -20'd95662}}, '{'{-20'd90089, 20'd15789, 20'd15789}, '{-20'd30649, -20'd118881, 20'd29720}, '{20'd29720, -20'd57583, -20'd74300}}, '{'{20'd6501, -20'd13003, -20'd90089}, '{-20'd22290, -20'd108664, -20'd88232}, '{-20'd75229, -20'd21361, -20'd53868}}, '{'{-20'd83588, -20'd72443, -20'd5573}, '{-20'd27863, -20'd53868, -20'd13931}, '{-20'd103092, -20'd20433, -20'd38079}}}
};
