localparam bit signed [0:10][15:0] Output4 = '{-16'd10315, -16'd16603, -16'd6998, -16'd11790, 16'd579, -16'd25215, -16'd7489, -16'd25462, -16'd16747, 16'd13576, -16'd7892};
