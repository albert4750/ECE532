localparam bit signed [0:2][0:31][0:4][0:4][24:0] Weight3 = '{
    '{'{'{25'd1955808, -25'd391162, 25'd2514611, 25'd111760, 25'd2794012}, '{-25'd335281, 25'd1452886, 25'd2179329, 25'd2291090, -25'd558802}, '{25'd2794012, 25'd1397006, 25'd4135138, 25'd3241054, 25'd111760}, '{25'd1508766, 25'd614683, 25'd391162, 25'd2123449, -25'd167641}, '{25'd1676407, 25'd111760, 25'd3408695, 25'd0, 25'd1955808}}, '{'{-25'd1899928, -25'd2682252, -25'd1508766, 25'd111760, 25'd1564647}, '{-25'd2402850, -25'd558802, -25'd1620527, -25'd782323, 25'd1732287}, '{-25'd1676407, -25'd391162, -25'd223521, 25'd1676407, 25'd949964}, '{-25'd279401, 25'd894084, -25'd838204, 25'd55880, 25'd1005844}, '{25'd2179329, 25'd2514611, -25'd782323, 25'd0, 25'd1899928}}, '{'{-25'd894084, 25'd1452886, 25'd2514611, 25'd2626371, 25'd894084}, '{25'd223521, -25'd223521, -25'd894084, -25'd1341126, -25'd223521}, '{25'd1229365, 25'd2235210, 25'd2011689, 25'd1899928, -25'd670563}, '{25'd0, -25'd1005844, 25'd1564647, 25'd1341126, 25'd1452886}, '{25'd502922, -25'd670563, 25'd2123449, -25'd1117605, -25'd502922}}, '{'{25'd614683, -25'd167641, 25'd1229365, 25'd1117605, -25'd111760}, '{25'd502922, 25'd614683, -25'd894084, -25'd1788168, 25'd335281}, '{-25'd1452886, 25'd1955808, 25'd1452886, -25'd447042, 25'd838204}, '{-25'd1229365, -25'd1564647, -25'd670563, 25'd1732287, 25'd1285246}, '{25'd335281, -25'd335281, -25'd782323, 25'd1117605, 25'd335281}}, '{'{-25'd447042, -25'd949964, -25'd1788168, -25'd838204, 25'd0}, '{25'd1397006, 25'd223521, -25'd614683, 25'd670563, 25'd447042}, '{-25'd670563, 25'd1732287, 25'd1564647, -25'd335281, 25'd502922}, '{25'd1117605, 25'd1285246, 25'd1397006, 25'd1173485, 25'd1229365}, '{-25'd670563, -25'd726443, 25'd1732287, 25'd55880, 25'd670563}}, '{'{25'd1061725, 25'd279401, -25'd726443, 25'd223521, -25'd223521}, '{-25'd1229365, -25'd1955808, -25'd782323, 25'd1173485, -25'd2179329}, '{-25'd391162, -25'd1508766, 25'd1508766, -25'd223521, 25'd614683}, '{-25'd1397006, -25'd1397006, 25'd1899928, -25'd279401, -25'd1899928}, '{25'd111760, -25'd558802, 25'd1620527, -25'd2179329, -25'd1341126}}, '{'{25'd614683, -25'd1061725, 25'd894084, -25'd1061725, 25'd1005844}, '{25'd726443, -25'd614683, -25'd1564647, 25'd1341126, -25'd670563}, '{25'd782323, 25'd502922, 25'd949964, 25'd335281, 25'd1117605}, '{-25'd391162, -25'd1005844, 25'd335281, -25'd1620527, -25'd2179329}, '{-25'd1564647, -25'd502922, 25'd1564647, -25'd111760, -25'd894084}}, '{'{-25'd1117605, -25'd2570491, 25'd2179329, -25'd279401, -25'd335281}, '{-25'd894084, -25'd2738132, 25'd1508766, 25'd279401, 25'd838204}, '{-25'd2235210, 25'd558802, 25'd3241054, 25'd2179329, -25'd335281}, '{-25'd2067569, -25'd1341126, -25'd502922, 25'd1676407, -25'd1620527}, '{-25'd1564647, -25'd3464575, 25'd614683, -25'd3352814, -25'd3017533}}, '{'{-25'd726443, -25'd223521, -25'd726443, -25'd1844048, 25'd167641}, '{-25'd391162, 25'd279401, 25'd279401, -25'd1341126, 25'd558802}, '{-25'd2570491, 25'd1788168, 25'd726443, 25'd2067569, 25'd1173485}, '{-25'd1341126, 25'd2067569, 25'd1173485, 25'd782323, -25'd447042}, '{-25'd2291090, 25'd335281, 25'd1508766, -25'd167641, -25'd447042}}, '{'{25'd4638060, -25'd782323, -25'd3129293, 25'd558802, 25'd5252743}, '{-25'd558802, -25'd4582180, -25'd5643904, 25'd502922, 25'd7096791}, '{25'd335281, -25'd3799856, -25'd6482108, -25'd949964, 25'd4805701}, '{25'd4861581, -25'd1173485, -25'd5308623, -25'd3632216, 25'd2514611}, '{25'd5923305, 25'd3520455, -25'd3632216, -25'd4749820, 25'd2291090}}, '{'{-25'd1620527, -25'd949964, -25'd335281, -25'd1117605, 25'd1229365}, '{-25'd1676407, -25'd894084, 25'd1229365, 25'd614683, -25'd670563}, '{25'd2067569, -25'd167641, 25'd838204, 25'd1117605, 25'd1676407}, '{25'd335281, 25'd670563, -25'd1452886, 25'd111760, 25'd0}, '{25'd949964, 25'd1117605, 25'd1397006, -25'd1620527, 25'd167641}}, '{'{-25'd894084, -25'd167641, -25'd614683, -25'd1452886, -25'd838204}, '{25'd1955808, 25'd1955808, -25'd447042, 25'd502922, -25'd1341126}, '{-25'd1005844, -25'd726443, 25'd1899928, -25'd1732287, -25'd502922}, '{-25'd726443, 25'd1732287, -25'd726443, 25'd502922, -25'd838204}, '{25'd1955808, 25'd502922, -25'd1285246, 25'd949964, -25'd670563}}, '{'{-25'd1788168, -25'd3352814, -25'd614683, -25'd335281, -25'd1899928}, '{-25'd1005844, -25'd3017533, 25'd1899928, -25'd949964, -25'd502922}, '{-25'd894084, 25'd949964, 25'd949964, 25'd3017533, 25'd782323}, '{25'd1117605, 25'd1117605, 25'd3799856, 25'd2067569, 25'd1452886}, '{-25'd1788168, -25'd3296934, -25'd1229365, -25'd1788168, 25'd335281}}, '{'{25'd279401, 25'd2011689, 25'd55880, -25'd167641, 25'd279401}, '{-25'd949964, -25'd1788168, -25'd1117605, 25'd1173485, -25'd614683}, '{-25'd726443, -25'd1564647, -25'd726443, -25'd447042, 25'd782323}, '{25'd670563, 25'd1564647, -25'd782323, 25'd223521, 25'd838204}, '{25'd670563, 25'd1508766, -25'd335281, -25'd1117605, -25'd1341126}}, '{'{25'd1620527, 25'd1452886, 25'd279401, 25'd1955808, 25'd111760}, '{25'd1564647, 25'd279401, 25'd502922, -25'd614683, -25'd670563}, '{25'd2011689, 25'd1676407, -25'd1564647, 25'd1173485, -25'd1061725}, '{-25'd1676407, -25'd1229365, 25'd1452886, 25'd1005844, 25'd614683}, '{-25'd1452886, 25'd2067569, 25'd447042, 25'd2011689, -25'd1005844}}, '{'{-25'd447042, 25'd838204, -25'd1341126, -25'd1117605, -25'd558802}, '{25'd447042, -25'd223521, -25'd1508766, -25'd726443, -25'd670563}, '{-25'd335281, -25'd279401, 25'd1061725, -25'd1005844, -25'd111760}, '{25'd1452886, 25'd1341126, -25'd614683, -25'd1732287, 25'd223521}, '{-25'd391162, 25'd949964, 25'd614683, -25'd726443, -25'd894084}}, '{'{25'd279401, -25'd1397006, -25'd167641, -25'd335281, -25'd1844048}, '{-25'd502922, 25'd1452886, 25'd167641, -25'd1620527, 25'd223521}, '{25'd2011689, 25'd502922, -25'd1732287, 25'd726443, 25'd1508766}, '{-25'd1285246, 25'd1229365, 25'd1452886, 25'd1620527, -25'd391162}, '{-25'd1788168, -25'd1676407, 25'd558802, 25'd111760, -25'd447042}}, '{'{25'd894084, -25'd1899928, -25'd894084, 25'd111760, -25'd1788168}, '{25'd1173485, 25'd894084, -25'd2179329, 25'd1452886, -25'd558802}, '{25'd894084, -25'd726443, 25'd949964, 25'd0, 25'd670563}, '{25'd502922, -25'd1955808, -25'd1564647, -25'd894084, -25'd1452886}, '{-25'd1117605, -25'd2067569, -25'd949964, -25'd1564647, -25'd1285246}}, '{'{25'd726443, -25'd2179329, -25'd279401, -25'd726443, -25'd558802}, '{25'd1620527, -25'd335281, -25'd1955808, -25'd838204, 25'd391162}, '{-25'd670563, 25'd1341126, -25'd558802, 25'd1285246, 25'd1620527}, '{-25'd223521, -25'd614683, 25'd782323, 25'd391162, -25'd2123449}, '{-25'd335281, -25'd1844048, -25'd1732287, -25'd782323, -25'd2067569}}, '{'{25'd1955808, 25'd1899928, 25'd1676407, -25'd167641, 25'd1117605}, '{-25'd670563, 25'd1005844, 25'd1452886, -25'd1564647, 25'd614683}, '{25'd1732287, -25'd1788168, -25'd223521, 25'd1005844, -25'd1452886}, '{25'd1285246, -25'd111760, -25'd279401, -25'd391162, -25'd55880}, '{-25'd726443, -25'd782323, -25'd1061725, 25'd335281, 25'd1117605}}, '{'{25'd2514611, 25'd3799856, 25'd4358659, 25'd3017533, -25'd1341126}, '{25'd167641, 25'd3911617, 25'd3352814, 25'd2626371, 25'd1397006}, '{25'd782323, 25'd4135138, 25'd5140982, 25'd614683, 25'd1452886}, '{-25'd1005844, 25'd111760, 25'd2682252, 25'd1844048, -25'd1732287}, '{-25'd2123449, -25'd335281, -25'd1899928, -25'd1285246, -25'd4358659}}, '{'{-25'd1508766, -25'd111760, 25'd1005844, -25'd1564647, 25'd502922}, '{25'd55880, 25'd1005844, -25'd1620527, -25'd1788168, 25'd1899928}, '{25'd0, 25'd1452886, 25'd223521, 25'd1955808, -25'd782323}, '{25'd55880, -25'd614683, 25'd1955808, -25'd55880, 25'd502922}, '{-25'd391162, 25'd1061725, 25'd1005844, -25'd1676407, 25'd949964}}, '{'{25'd726443, 25'd1788168, 25'd1341126, 25'd614683, -25'd223521}, '{25'd0, -25'd838204, 25'd3129293, 25'd223521, 25'd2738132}, '{-25'd1285246, 25'd2011689, 25'd1229365, 25'd558802, 25'd1508766}, '{25'd2067569, 25'd335281, 25'd3129293, 25'd167641, -25'd558802}, '{-25'd894084, 25'd2682252, -25'd279401, 25'd1676407, 25'd1899928}}, '{'{-25'd782323, -25'd2067569, 25'd558802, 25'd1061725, -25'd1061725}, '{-25'd55880, -25'd1341126, 25'd1117605, -25'd1788168, 25'd1173485}, '{25'd614683, -25'd1620527, -25'd1005844, 25'd614683, 25'd949964}, '{-25'd2067569, -25'd167641, 25'd726443, -25'd1620527, 25'd2235210}, '{-25'd167641, 25'd223521, -25'd2291090, 25'd1397006, 25'd2179329}}, '{'{25'd1452886, -25'd335281, -25'd838204, 25'd782323, 25'd1676407}, '{25'd670563, -25'd1117605, 25'd1564647, -25'd1117605, 25'd1620527}, '{-25'd279401, -25'd1620527, -25'd838204, 25'd167641, -25'd782323}, '{25'd1732287, -25'd55880, 25'd1005844, -25'd558802, -25'd894084}, '{-25'd279401, 25'd1229365, -25'd558802, -25'd1117605, -25'd670563}}, '{'{25'd894084, -25'd838204, -25'd1564647, -25'd1955808, -25'd3017533}, '{25'd111760, -25'd167641, 25'd223521, -25'd1341126, -25'd2346970}, '{-25'd1173485, -25'd1676407, -25'd1452886, -25'd2849892, 25'd1005844}, '{-25'd670563, -25'd2179329, -25'd838204, 25'd391162, -25'd391162}, '{-25'd2123449, -25'd223521, -25'd2794012, 25'd670563, -25'd447042}}, '{'{-25'd1061725, 25'd1508766, -25'd391162, 25'd1229365, -25'd335281}, '{-25'd1005844, 25'd782323, -25'd670563, -25'd1173485, -25'd2123449}, '{-25'd558802, 25'd2570491, 25'd391162, 25'd894084, -25'd447042}, '{-25'd1117605, 25'd1397006, 25'd838204, -25'd838204, -25'd167641}, '{-25'd502922, -25'd670563, 25'd335281, -25'd2402850, -25'd55880}}, '{'{25'd1452886, 25'd670563, -25'd447042, 25'd894084, 25'd1844048}, '{-25'd558802, 25'd1285246, 25'd726443, 25'd502922, -25'd335281}, '{-25'd670563, -25'd1341126, -25'd391162, -25'd782323, -25'd447042}, '{25'd167641, 25'd1397006, 25'd1005844, -25'd167641, 25'd726443}, '{25'd1397006, 25'd1564647, 25'd335281, -25'd1508766, -25'd55880}}, '{'{25'd1676407, -25'd1061725, -25'd335281, 25'd670563, -25'd1173485}, '{-25'd1732287, 25'd1397006, -25'd838204, 25'd1732287, 25'd838204}, '{-25'd1341126, -25'd1564647, 25'd279401, 25'd726443, -25'd614683}, '{25'd949964, -25'd1508766, -25'd1732287, 25'd1955808, 25'd1899928}, '{25'd1899928, -25'd726443, 25'd1285246, 25'd1397006, -25'd279401}}, '{'{-25'd1844048, 25'd167641, 25'd223521, -25'd1341126, -25'd1341126}, '{-25'd502922, -25'd335281, 25'd1620527, 25'd949964, 25'd670563}, '{25'd782323, 25'd1676407, 25'd1173485, 25'd670563, 25'd2067569}, '{-25'd558802, 25'd1564647, -25'd614683, 25'd726443, -25'd838204}, '{25'd1955808, 25'd670563, 25'd1117605, 25'd502922, -25'd726443}}, '{'{-25'd838204, 25'd1229365, -25'd55880, 25'd1117605, -25'd894084}, '{25'd1676407, -25'd894084, -25'd1676407, 25'd949964, -25'd223521}, '{-25'd558802, 25'd1173485, 25'd1173485, 25'd838204, 25'd279401}, '{25'd55880, 25'd1285246, -25'd1341126, -25'd502922, 25'd949964}, '{25'd670563, 25'd335281, -25'd1173485, 25'd782323, 25'd0}}, '{'{25'd1285246, 25'd894084, -25'd1229365, -25'd447042, 25'd1229365}, '{25'd1564647, 25'd2067569, -25'd1061725, 25'd949964, 25'd335281}, '{-25'd1676407, -25'd1620527, -25'd1341126, -25'd111760, -25'd782323}, '{25'd2067569, 25'd1732287, -25'd502922, -25'd55880, 25'd1899928}, '{25'd1005844, -25'd949964, -25'd1397006, 25'd1173485, 25'd2011689}}},
    '{'{'{25'd0, -25'd2969436, 25'd379077, 25'd1263590, -25'd1769026}, '{-25'd1200410, -25'd1642667, -25'd821333, 25'd505436, 25'd315897}, '{25'd1705846, -25'd947692, -25'd1074051, -25'd1453128, -25'd126359}, '{25'd631795, 25'd126359, -25'd1705846, -25'd884513, -25'd2274462}, '{-25'd2274462, -25'd1453128, -25'd2464000, -25'd1200410, -25'd1137231}}, '{'{-25'd189538, -25'd758154, -25'd758154, -25'd694974, 25'd694974}, '{-25'd2148103, -25'd63179, -25'd694974, 25'd315897, 25'd2148103}, '{25'd379077, 25'd0, -25'd1958564, 25'd315897, 25'd947692}, '{-25'd1579487, -25'd63179, -25'd2084923, -25'd568615, 25'd1832205}, '{-25'd1705846, 25'd252718, 25'd884513, 25'd442256, 25'd631795}}, '{'{-25'd442256, -25'd1895385, -25'd758154, -25'd947692, -25'd2021744}, '{25'd0, 25'd758154, -25'd884513, -25'd568615, -25'd1705846}, '{25'd694974, -25'd1326769, 25'd568615, -25'd379077, -25'd821333}, '{-25'd1074051, 25'd1074051, 25'd758154, 25'd189538, 25'd126359}, '{25'd1453128, -25'd2021744, 25'd568615, 25'd189538, -25'd1579487}}, '{'{25'd1200410, -25'd1579487, 25'd379077, 25'd1389949, 25'd1200410}, '{25'd126359, 25'd1705846, -25'd1389949, 25'd884513, 25'd189538}, '{-25'd1326769, 25'd1832205, -25'd1326769, -25'd1137231, 25'd631795}, '{-25'd947692, 25'd2084923, -25'd1769026, -25'd947692, 25'd821333}, '{25'd1074051, -25'd884513, 25'd821333, -25'd947692, -25'd1137231}}, '{'{25'd568615, -25'd758154, 25'd1958564, -25'd1263590, -25'd505436}, '{25'd758154, 25'd2021744, 25'd505436, 25'd1579487, 25'd2084923}, '{25'd947692, 25'd1389949, -25'd252718, -25'd1137231, 25'd1010872}, '{-25'd1453128, 25'd821333, 25'd126359, 25'd189538, 25'd1895385}, '{-25'd505436, 25'd1200410, -25'd1137231, 25'd2148103, 25'd1958564}}, '{'{-25'd1200410, -25'd1326769, -25'd821333, -25'd1074051, -25'd505436}, '{-25'd1642667, 25'd694974, -25'd252718, 25'd1769026, -25'd1010872}, '{-25'd1832205, 25'd126359, -25'd1074051, 25'd821333, -25'd631795}, '{-25'd2021744, 25'd252718, 25'd315897, -25'd2021744, -25'd252718}, '{-25'd1516308, 25'd884513, -25'd1769026, 25'd379077, -25'd1200410}}, '{'{25'd315897, 25'd0, 25'd1453128, -25'd631795, 25'd821333}, '{25'd1453128, 25'd379077, 25'd1389949, -25'd315897, -25'd694974}, '{25'd884513, 25'd126359, -25'd1074051, 25'd1074051, -25'd758154}, '{-25'd1516308, -25'd189538, -25'd821333, 25'd1010872, -25'd315897}, '{-25'd694974, 25'd758154, -25'd947692, -25'd884513, 25'd1389949}}, '{'{-25'd1705846, 25'd631795, 25'd1453128, -25'd821333, 25'd442256}, '{-25'd694974, 25'd379077, 25'd1326769, -25'd1389949, 25'd315897}, '{25'd631795, -25'd568615, 25'd2653539, 25'd1832205, -25'd379077}, '{25'd63179, -25'd3032616, 25'd252718, -25'd1137231, 25'd884513}, '{-25'd3158975, -25'd505436, -25'd1705846, -25'd3474872, -25'd758154}}, '{'{-25'd2464000, -25'd2590359, -25'd1200410, -25'd884513, -25'd1263590}, '{-25'd1958564, -25'd3095795, -25'd505436, 25'd947692, -25'd1074051}, '{25'd694974, 25'd1137231, 25'd442256, -25'd1769026, 25'd568615}, '{-25'd1958564, -25'd1010872, 25'd2464000, -25'd1453128, 25'd315897}, '{-25'd379077, 25'd1137231, 25'd2021744, -25'd2211282, 25'd694974}}, '{'{25'd1642667, -25'd379077, -25'd1453128, -25'd1579487, 25'd5749334}, '{-25'd1769026, -25'd2211282, -25'd4801641, -25'd1705846, 25'd6317949}, '{25'd2400821, -25'd442256, -25'd6128411, -25'd4485744, 25'd7202462}, '{25'd2021744, 25'd1074051, -25'd4485744, -25'd4928000, 25'd189538}, '{25'd8023796, 25'd6191590, -25'd442256, -25'd2716718, -25'd505436}}, '{'{25'd505436, 25'd2148103, -25'd505436, -25'd189538, -25'd315897}, '{25'd2021744, 25'd1895385, -25'd252718, -25'd758154, 25'd379077}, '{-25'd947692, -25'd884513, -25'd568615, -25'd1137231, 25'd1137231}, '{25'd442256, 25'd1453128, 25'd1389949, -25'd379077, -25'd379077}, '{-25'd821333, 25'd1200410, -25'd568615, -25'd758154, 25'd884513}}, '{'{25'd2148103, -25'd1137231, 25'd1389949, -25'd1263590, 25'd568615}, '{-25'd1263590, -25'd189538, 25'd1579487, 25'd2148103, -25'd315897}, '{25'd631795, 25'd442256, -25'd1579487, 25'd1074051, 25'd1263590}, '{-25'd189538, -25'd252718, -25'd694974, 25'd1705846, 25'd694974}, '{25'd1769026, 25'd2084923, -25'd442256, 25'd1832205, -25'd1389949}}, '{'{25'd1200410, -25'd1895385, -25'd631795, -25'd126359, -25'd1074051}, '{-25'd2400821, -25'd2274462, 25'd63179, 25'd189538, -25'd2148103}, '{25'd1010872, -25'd2464000, 25'd3980308, 25'd442256, 25'd0}, '{-25'd252718, -25'd2906257, 25'd1074051, -25'd1200410, -25'd1579487}, '{25'd1705846, 25'd126359, -25'd126359, 25'd126359, -25'd1895385}}, '{'{25'd1832205, -25'd1389949, 25'd1453128, -25'd1074051, -25'd1074051}, '{25'd1263590, -25'd758154, 25'd442256, -25'd758154, -25'd1263590}, '{25'd1074051, -25'd315897, 25'd2021744, 25'd1895385, 25'd1516308}, '{25'd0, -25'd379077, 25'd63179, -25'd694974, -25'd1579487}, '{25'd1010872, 25'd1010872, 25'd1074051, -25'd1137231, -25'd821333}}, '{'{25'd442256, 25'd1326769, -25'd1769026, -25'd1200410, -25'd947692}, '{25'd126359, -25'd189538, 25'd189538, 25'd1200410, -25'd1895385}, '{-25'd1010872, -25'd252718, -25'd1453128, 25'd1579487, -25'd1705846}, '{-25'd442256, 25'd1958564, -25'd631795, 25'd315897, 25'd1705846}, '{25'd1263590, -25'd947692, -25'd1453128, 25'd505436, 25'd568615}}, '{'{-25'd1137231, 25'd2274462, -25'd1263590, -25'd1516308, -25'd315897}, '{-25'd1074051, 25'd63179, 25'd1200410, -25'd1137231, 25'd1958564}, '{-25'd63179, 25'd2148103, 25'd2653539, 25'd568615, -25'd884513}, '{-25'd1769026, 25'd2148103, -25'd189538, 25'd694974, 25'd0}, '{25'd1579487, -25'd947692, -25'd821333, -25'd1263590, -25'd631795}}, '{'{-25'd63179, 25'd1453128, -25'd1074051, 25'd1832205, 25'd1200410}, '{-25'd694974, -25'd315897, -25'd315897, -25'd1453128, -25'd758154}, '{-25'd1010872, 25'd1074051, 25'd1389949, 25'd1958564, 25'd884513}, '{25'd315897, 25'd1200410, 25'd1516308, 25'd694974, 25'd884513}, '{-25'd1137231, -25'd1705846, 25'd315897, -25'd884513, 25'd1642667}}, '{'{-25'd505436, -25'd1832205, 25'd189538, -25'd694974, -25'd631795}, '{-25'd884513, 25'd758154, 25'd2021744, 25'd568615, 25'd126359}, '{-25'd1579487, -25'd1200410, -25'd1579487, 25'd1010872, 25'd1074051}, '{25'd1263590, -25'd505436, 25'd63179, 25'd821333, -25'd1769026}, '{25'd442256, -25'd1074051, -25'd1705846, 25'd1137231, -25'd1769026}}, '{'{-25'd1389949, 25'd631795, 25'd884513, 25'd694974, 25'd379077}, '{25'd1895385, 25'd884513, 25'd379077, 25'd1263590, 25'd189538}, '{-25'd1516308, 25'd947692, 25'd2021744, 25'd315897, 25'd189538}, '{25'd379077, 25'd1832205, 25'd1326769, 25'd63179, -25'd1200410}, '{25'd1642667, -25'd1705846, 25'd1769026, 25'd126359, -25'd1263590}}, '{'{25'd315897, 25'd189538, 25'd1958564, -25'd126359, 25'd1769026}, '{25'd126359, 25'd1389949, 25'd442256, -25'd63179, 25'd568615}, '{-25'd1453128, 25'd1769026, 25'd1453128, 25'd505436, 25'd1074051}, '{-25'd315897, -25'd1642667, 25'd1832205, 25'd1453128, 25'd1010872}, '{25'd1137231, 25'd1958564, 25'd631795, -25'd568615, -25'd1705846}}, '{'{25'd3601231, 25'd3601231, 25'd5559795, 25'd4043488, 25'd2211282}, '{25'd2211282, 25'd4169847, 25'd4991180, 25'd5559795, 25'd1263590}, '{25'd2400821, 25'd4359385, 25'd6317949, 25'd4043488, 25'd2084923}, '{25'd315897, 25'd2716718, 25'd2779898, 25'd3285334, 25'd694974}, '{25'd252718, 25'd1453128, 25'd1010872, 25'd758154, -25'd694974}}, '{'{-25'd884513, 25'd505436, 25'd442256, 25'd947692, -25'd1263590}, '{25'd1010872, 25'd821333, -25'd694974, 25'd2400821, 25'd379077}, '{25'd947692, 25'd126359, -25'd315897, 25'd1453128, 25'd694974}, '{25'd1895385, -25'd1074051, 25'd821333, -25'd884513, 25'd1074051}, '{-25'd1200410, 25'd189538, 25'd1010872, -25'd379077, 25'd568615}}, '{'{-25'd2211282, -25'd821333, 25'd2021744, 25'd442256, 25'd252718}, '{-25'd2590359, -25'd1074051, -25'd884513, 25'd884513, 25'd568615}, '{-25'd2211282, 25'd821333, -25'd821333, 25'd63179, -25'd126359}, '{25'd947692, 25'd1389949, 25'd631795, 25'd189538, -25'd884513}, '{25'd189538, -25'd1263590, 25'd1200410, -25'd1895385, -25'd1074051}}, '{'{25'd1895385, 25'd2274462, -25'd821333, -25'd2084923, -25'd947692}, '{25'd947692, 25'd1895385, -25'd2021744, 25'd694974, 25'd1958564}, '{25'd2527180, 25'd568615, -25'd1389949, -25'd2084923, -25'd821333}, '{25'd2906257, -25'd884513, 25'd189538, -25'd379077, -25'd947692}, '{25'd1137231, 25'd0, -25'd884513, -25'd2906257, 25'd1200410}}, '{'{25'd1832205, 25'd1389949, -25'd1579487, -25'd1769026, 25'd694974}, '{25'd821333, 25'd63179, -25'd1642667, 25'd442256, 25'd1263590}, '{-25'd758154, -25'd568615, -25'd1326769, -25'd442256, -25'd884513}, '{25'd758154, 25'd315897, 25'd1389949, 25'd1705846, 25'd1705846}, '{25'd1200410, -25'd568615, 25'd505436, -25'd1200410, -25'd1389949}}, '{'{25'd694974, 25'd694974, -25'd631795, -25'd947692, -25'd1895385}, '{-25'd758154, -25'd1200410, -25'd2779898, -25'd2400821, -25'd1453128}, '{-25'd252718, -25'd505436, -25'd2653539, -25'd2653539, 25'd379077}, '{-25'd63179, -25'd694974, -25'd1010872, -25'd1895385, -25'd1832205}, '{-25'd442256, 25'd189538, 25'd0, -25'd947692, -25'd1389949}}, '{'{-25'd2653539, 25'd1010872, -25'd1326769, 25'd1389949, -25'd63179}, '{-25'd63179, -25'd1705846, 25'd1263590, 25'd568615, -25'd1958564}, '{-25'd1074051, 25'd1389949, 25'd1642667, 25'd2021744, -25'd1579487}, '{-25'd694974, 25'd821333, -25'd1074051, -25'd1516308, -25'd1010872}, '{-25'd2021744, -25'd1263590, -25'd1389949, 25'd2464000, -25'd379077}}, '{'{25'd189538, -25'd252718, -25'd1389949, 25'd1769026, -25'd252718}, '{-25'd1705846, 25'd1642667, -25'd252718, -25'd1137231, 25'd1516308}, '{25'd1200410, 25'd1642667, 25'd442256, -25'd568615, -25'd1769026}, '{-25'd1769026, -25'd1074051, -25'd1769026, 25'd63179, -25'd126359}, '{-25'd1389949, 25'd1200410, 25'd1389949, -25'd379077, -25'd252718}}, '{'{-25'd63179, 25'd189538, 25'd884513, 25'd821333, -25'd1137231}, '{25'd1958564, 25'd63179, -25'd63179, 25'd0, 25'd1895385}, '{25'd947692, 25'd758154, 25'd1137231, -25'd631795, -25'd505436}, '{25'd2021744, -25'd63179, -25'd568615, -25'd1453128, -25'd568615}, '{25'd568615, 25'd1263590, 25'd505436, 25'd1263590, -25'd1010872}}, '{'{-25'd1705846, 25'd947692, -25'd947692, 25'd2021744, -25'd694974}, '{25'd252718, 25'd442256, 25'd821333, -25'd821333, -25'd1705846}, '{25'd1769026, 25'd1769026, -25'd505436, -25'd1137231, 25'd1453128}, '{25'd758154, 25'd1642667, 25'd884513, 25'd1010872, -25'd1010872}, '{-25'd758154, 25'd1516308, 25'd1958564, -25'd1389949, -25'd379077}}, '{'{-25'd505436, 25'd631795, -25'd568615, -25'd1579487, -25'd694974}, '{-25'd821333, -25'd1705846, 25'd694974, -25'd1263590, -25'd442256}, '{-25'd189538, -25'd505436, 25'd1579487, 25'd1958564, 25'd568615}, '{-25'd315897, 25'd442256, -25'd1705846, -25'd884513, 25'd568615}, '{25'd1516308, 25'd0, -25'd694974, -25'd1579487, 25'd694974}}, '{'{-25'd442256, 25'd252718, 25'd1832205, 25'd1389949, 25'd1705846}, '{25'd1453128, -25'd315897, 25'd1200410, 25'd568615, 25'd2084923}, '{-25'd884513, 25'd1389949, 25'd1895385, -25'd758154, -25'd821333}, '{25'd1705846, -25'd694974, 25'd1137231, -25'd1200410, -25'd1579487}, '{-25'd884513, -25'd1326769, -25'd821333, 25'd1705846, 25'd821333}}},
    '{'{'{-25'd1245793, 25'd0, 25'd389310, -25'd77862, -25'd233586}, '{-25'd2803035, -25'd1323655, -25'd856483, -25'd545035, -25'd2180138}, '{-25'd1012207, -25'd1090069, -25'd622897, 25'd389310, 25'd233586}, '{-25'd2024414, 25'd77862, -25'd1868690, -25'd700759, -25'd1790828}, '{-25'd3659518, -25'd3348070, -25'd233586, -25'd2880897, -25'd1245793}}, '{'{25'd155724, 25'd1323655, -25'd545035, 25'd1167931, 25'd545035}, '{25'd1479380, -25'd155724, 25'd0, 25'd622897, -25'd233586}, '{-25'd467173, 25'd467173, -25'd1790828, -25'd311448, -25'd934345}, '{25'd2335863, -25'd389310, -25'd1401518, -25'd1635104, 25'd1401518}, '{25'd1712966, -25'd1557242, 25'd467173, 25'd1090069, 25'd1167931}}, '{'{-25'd1090069, -25'd1323655, 25'd1790828, -25'd1401518, -25'd856483}, '{-25'd1245793, -25'd1790828, 25'd233586, -25'd856483, -25'd1790828}, '{-25'd311448, 25'd1090069, -25'd778621, -25'd1479380, -25'd1323655}, '{-25'd77862, -25'd1479380, 25'd778621, 25'd389310, 25'd1012207}, '{25'd77862, 25'd934345, -25'd155724, -25'd1635104, 25'd1635104}}, '{'{25'd467173, 25'd0, 25'd1635104, 25'd1712966, -25'd1167931}, '{25'd1557242, 25'd233586, 25'd1712966, 25'd2102276, -25'd1479380}, '{25'd0, -25'd77862, -25'd311448, 25'd856483, -25'd856483}, '{25'd622897, 25'd233586, -25'd545035, -25'd233586, -25'd1635104}, '{25'd1323655, 25'd1012207, -25'd1557242, 25'd1868690, 25'd1712966}}, '{'{-25'd856483, 25'd311448, 25'd1557242, 25'd622897, 25'd0}, '{25'd311448, -25'd1401518, 25'd2180138, 25'd311448, 25'd1167931}, '{25'd700759, 25'd1401518, -25'd1479380, 25'd700759, -25'd389310}, '{-25'd1245793, -25'd1712966, -25'd622897, 25'd1557242, -25'd1401518}, '{-25'd389310, -25'd1012207, -25'd1245793, 25'd2180138, 25'd1090069}}, '{'{25'd934345, -25'd389310, 25'd700759, -25'd622897, -25'd311448}, '{-25'd1012207, -25'd1323655, 25'd2180138, 25'd1479380, 25'd1790828}, '{-25'd233586, -25'd934345, 25'd2258001, 25'd311448, -25'd1946552}, '{25'd1635104, -25'd155724, 25'd1712966, 25'd233586, 25'd233586}, '{25'd1012207, 25'd1323655, 25'd1012207, -25'd1090069, -25'd155724}}, '{'{25'd1946552, 25'd1868690, -25'd1167931, -25'd77862, 25'd856483}, '{-25'd233586, -25'd1323655, 25'd233586, 25'd77862, 25'd934345}, '{25'd1557242, 25'd545035, 25'd2258001, 25'd77862, -25'd389310}, '{-25'd1090069, 25'd934345, -25'd700759, 25'd778621, 25'd622897}, '{-25'd1245793, 25'd622897, 25'd778621, -25'd1868690, 25'd2102276}}, '{'{-25'd700759, 25'd1167931, 25'd2803035, 25'd2880897, 25'd1323655}, '{25'd77862, 25'd3270208, 25'd5761794, 25'd2180138, 25'd1557242}, '{25'd4048829, 25'd3893104, 25'd5061036, 25'd3737380, 25'd2258001}, '{25'd0, 25'd3737380, 25'd5216760, 25'd3659518, 25'd1401518}, '{-25'd934345, 25'd1557242, 25'd856483, 25'd778621, -25'd622897}}, '{'{-25'd1790828, -25'd233586, -25'd155724, 25'd622897, -25'd1946552}, '{-25'd2413725, -25'd1012207, -25'd1790828, 25'd1090069, 25'd77862}, '{25'd155724, 25'd1557242, -25'd155724, 25'd467173, -25'd1479380}, '{-25'd1790828, 25'd1323655, 25'd934345, -25'd1635104, -25'd545035}, '{-25'd934345, 25'd2102276, 25'd934345, 25'd155724, 25'd545035}}, '{'{-25'd77862, -25'd3036621, -25'd4671725, -25'd1635104, 25'd8798416}, '{-25'd3348070, -25'd6851864, -25'd5294622, -25'd389310, 25'd6151105}, '{25'd2803035, -25'd2880897, -25'd2725173, -25'd1167931, 25'd8798416}, '{25'd4905311, 25'd1090069, -25'd4282415, -25'd2880897, 25'd1323655}, '{25'd9888485, 25'd8564830, 25'd77862, -25'd2180138, 25'd389310}}, '{'{25'd0, -25'd545035, -25'd311448, 25'd778621, 25'd622897}, '{25'd0, 25'd1245793, -25'd700759, 25'd622897, 25'd545035}, '{-25'd389310, 25'd1479380, 25'd1401518, 25'd700759, 25'd622897}, '{25'd1245793, 25'd1401518, -25'd1401518, -25'd1557242, 25'd934345}, '{25'd1479380, -25'd1557242, -25'd1635104, 25'd1245793, 25'd1557242}}, '{'{-25'd155724, 25'd1401518, -25'd467173, -25'd1012207, -25'd1090069}, '{-25'd1479380, 25'd1635104, -25'd622897, 25'd1401518, 25'd856483}, '{25'd311448, 25'd2024414, 25'd1557242, -25'd389310, 25'd1090069}, '{25'd1323655, 25'd856483, -25'd856483, 25'd856483, -25'd1245793}, '{25'd2258001, 25'd934345, -25'd155724, -25'd934345, -25'd545035}}, '{'{-25'd1245793, -25'd2647311, 25'd1868690, -25'd1946552, 25'd934345}, '{-25'd2803035, -25'd2024414, -25'd700759, -25'd1167931, -25'd3503794}, '{25'd1712966, -25'd1946552, 25'd3036621, 25'd778621, -25'd389310}, '{-25'd934345, -25'd1245793, -25'd1635104, -25'd2880897, -25'd934345}, '{25'd700759, -25'd1479380, 25'd1167931, 25'd77862, -25'd1012207}}, '{'{-25'd778621, 25'd155724, -25'd700759, 25'd467173, 25'd1401518}, '{25'd1868690, -25'd1090069, -25'd1012207, 25'd1323655, -25'd77862}, '{-25'd700759, 25'd0, 25'd2102276, 25'd2102276, 25'd1323655}, '{-25'd233586, -25'd1401518, 25'd622897, -25'd1712966, 25'd1868690}, '{-25'd1790828, 25'd1557242, -25'd1323655, -25'd856483, -25'd1712966}}, '{'{-25'd77862, 25'd934345, 25'd934345, -25'd1012207, 25'd1712966}, '{25'd1946552, -25'd1323655, -25'd389310, -25'd1012207, 25'd1712966}, '{-25'd233586, -25'd1557242, 25'd77862, -25'd155724, -25'd233586}, '{-25'd77862, 25'd2258001, -25'd622897, 25'd1946552, 25'd856483}, '{25'd934345, 25'd1012207, 25'd1635104, 25'd2024414, -25'd545035}}, '{'{-25'd155724, 25'd233586, 25'd2024414, -25'd778621, -25'd2024414}, '{25'd1946552, 25'd2491587, 25'd1790828, 25'd1712966, -25'd467173}, '{25'd1790828, 25'd1401518, -25'd1401518, -25'd2102276, -25'd77862}, '{25'd1090069, 25'd311448, -25'd856483, 25'd1401518, -25'd2258001}, '{-25'd311448, -25'd1635104, -25'd1401518, 25'd700759, -25'd622897}}, '{'{25'd1790828, -25'd1479380, -25'd467173, -25'd155724, -25'd1167931}, '{25'd856483, 25'd1401518, -25'd1401518, -25'd467173, -25'd1167931}, '{25'd311448, 25'd856483, 25'd934345, -25'd77862, -25'd1245793}, '{25'd155724, 25'd311448, -25'd545035, 25'd1401518, 25'd2102276}, '{-25'd856483, -25'd856483, 25'd1401518, -25'd1790828, 25'd545035}}, '{'{-25'd1790828, -25'd1012207, -25'd1090069, -25'd1245793, -25'd1090069}, '{-25'd1712966, 25'd545035, 25'd1323655, 25'd233586, 25'd856483}, '{25'd77862, 25'd77862, 25'd1790828, -25'd1479380, 25'd778621}, '{-25'd1323655, 25'd233586, 25'd389310, 25'd1790828, 25'd1167931}, '{25'd1245793, -25'd1868690, -25'd934345, 25'd1323655, 25'd856483}}, '{'{-25'd311448, -25'd622897, 25'd0, 25'd545035, -25'd2102276}, '{25'd1167931, 25'd1323655, 25'd2024414, 25'd856483, -25'd1245793}, '{25'd934345, -25'd1090069, 25'd1635104, -25'd622897, 25'd77862}, '{-25'd1790828, -25'd1868690, -25'd467173, 25'd1557242, -25'd622897}, '{-25'd233586, -25'd155724, -25'd622897, -25'd934345, 25'd778621}}, '{'{-25'd1401518, 25'd934345, -25'd1323655, 25'd622897, -25'd1323655}, '{25'd1479380, 25'd1090069, -25'd622897, 25'd2024414, 25'd233586}, '{-25'd1479380, -25'd1167931, 25'd856483, -25'd1635104, -25'd233586}, '{25'd934345, 25'd1635104, -25'd1012207, 25'd467173, 25'd1635104}, '{-25'd934345, -25'd77862, -25'd545035, -25'd467173, -25'd77862}}, '{'{25'd545035, 25'd2803035, 25'd3114483, 25'd311448, 25'd934345}, '{25'd2725173, 25'd4282415, 25'd2880897, 25'd1712966, -25'd1245793}, '{25'd1946552, 25'd1557242, 25'd3893104, 25'd545035, 25'd2102276}, '{-25'd1323655, -25'd155724, -25'd311448, -25'd1712966, -25'd2258001}, '{-25'd622897, 25'd77862, 25'd622897, -25'd1790828, -25'd3893104}}, '{'{-25'd1012207, 25'd934345, -25'd622897, 25'd1479380, -25'd389310}, '{-25'd622897, 25'd1557242, -25'd77862, 25'd1167931, -25'd1790828}, '{25'd1635104, -25'd1712966, 25'd1479380, 25'd77862, -25'd700759}, '{-25'd1012207, 25'd856483, -25'd1323655, -25'd1635104, 25'd778621}, '{-25'd1946552, 25'd700759, -25'd545035, -25'd1868690, -25'd545035}}, '{'{-25'd934345, -25'd3581656, -25'd389310, -25'd311448, -25'd77862}, '{-25'd2569449, -25'd1245793, -25'd2102276, -25'd1790828, -25'd389310}, '{-25'd3192346, -25'd155724, -25'd3114483, -25'd389310, -25'd3270208}, '{-25'd3737380, -25'd2335863, -25'd1790828, -25'd1245793, -25'd77862}, '{-25'd3036621, -25'd1012207, -25'd155724, -25'd1790828, -25'd3114483}}, '{'{25'd389310, 25'd622897, -25'd1401518, -25'd1868690, 25'd856483}, '{25'd545035, -25'd622897, 25'd0, 25'd467173, 25'd934345}, '{-25'd155724, 25'd1323655, -25'd1401518, 25'd1401518, 25'd77862}, '{25'd700759, -25'd856483, -25'd1012207, -25'd1479380, 25'd1479380}, '{25'd1245793, 25'd1557242, -25'd1712966, -25'd77862, 25'd1868690}}, '{'{25'd1167931, 25'd1012207, -25'd311448, -25'd778621, -25'd778621}, '{25'd389310, 25'd467173, 25'd389310, 25'd856483, 25'd934345}, '{-25'd934345, 25'd155724, 25'd1946552, 25'd1635104, 25'd2102276}, '{-25'd1557242, -25'd1012207, 25'd1090069, 25'd1090069, 25'd1635104}, '{-25'd1557242, 25'd1557242, -25'd1090069, 25'd1790828, 25'd1868690}}, '{'{-25'd155724, -25'd1090069, 25'd467173, -25'd3036621, 25'd778621}, '{25'd389310, -25'd2569449, 25'd0, 25'd934345, -25'd2725173}, '{-25'd2647311, -25'd2024414, -25'd2569449, 25'd700759, -25'd1635104}, '{-25'd2335863, -25'd77862, -25'd1012207, 25'd0, -25'd2958759}, '{-25'd1090069, -25'd545035, 25'd233586, 25'd934345, 25'd700759}}, '{'{25'd0, 25'd3581656, 25'd1790828, 25'd0, 25'd2958759}, '{25'd1245793, 25'd545035, 25'd3581656, 25'd2958759, 25'd1323655}, '{-25'd2491587, 25'd389310, -25'd1245793, -25'd934345, -25'd1245793}, '{-25'd1790828, -25'd1868690, 25'd1401518, 25'd778621, 25'd1090069}, '{-25'd2102276, -25'd1712966, -25'd622897, 25'd545035, 25'd77862}}, '{'{25'd2102276, 25'd1090069, 25'd934345, -25'd77862, -25'd1557242}, '{-25'd1401518, -25'd1401518, -25'd1635104, 25'd311448, 25'd1946552}, '{25'd1946552, 25'd2258001, 25'd856483, 25'd1557242, 25'd1946552}, '{25'd1245793, -25'd1012207, 25'd700759, -25'd233586, -25'd1635104}, '{-25'd856483, 25'd77862, 25'd1868690, 25'd1557242, 25'd389310}}, '{'{25'd934345, -25'd622897, -25'd389310, 25'd1479380, -25'd934345}, '{25'd1323655, 25'd311448, -25'd622897, -25'd311448, 25'd1245793}, '{-25'd1012207, -25'd311448, -25'd1712966, -25'd1635104, 25'd1557242}, '{25'd2180138, -25'd700759, -25'd1712966, 25'd1090069, 25'd155724}, '{25'd1557242, 25'd1479380, -25'd545035, -25'd934345, 25'd77862}}, '{'{25'd856483, -25'd1635104, 25'd545035, 25'd2024414, -25'd1167931}, '{25'd311448, -25'd1401518, -25'd545035, -25'd1167931, -25'd77862}, '{25'd1323655, 25'd545035, -25'd1323655, -25'd1479380, 25'd1946552}, '{-25'd1323655, -25'd700759, 25'd622897, 25'd0, -25'd934345}, '{25'd233586, -25'd934345, 25'd1012207, -25'd233586, 25'd856483}}, '{'{25'd2335863, -25'd1479380, 25'd2102276, 25'd389310, -25'd1557242}, '{25'd311448, 25'd856483, -25'd233586, 25'd389310, 25'd1712966}, '{-25'd467173, 25'd467173, -25'd622897, 25'd389310, 25'd467173}, '{-25'd778621, -25'd155724, 25'd1712966, -25'd467173, 25'd1167931}, '{-25'd1323655, 25'd1479380, 25'd856483, 25'd2102276, -25'd778621}}, '{'{25'd856483, -25'd1401518, -25'd233586, 25'd1712966, -25'd467173}, '{25'd233586, 25'd1635104, 25'd700759, 25'd1946552, 25'd155724}, '{25'd2024414, 25'd700759, -25'd233586, 25'd467173, -25'd389310}, '{-25'd856483, 25'd2180138, 25'd1790828, -25'd934345, -25'd311448}, '{25'd778621, -25'd1245793, -25'd545035, -25'd1245793, 25'd1479380}}}
};
