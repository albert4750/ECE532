localparam bit signed [0:2][47:0] Bias3 = '{-48'd72278, -48'd44950, -48'd4483};
