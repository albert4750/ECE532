localparam bit signed [0:26][19:0] Output5 = '{-20'd92, 20'd58, -20'd179, -20'd87, 20'd91, -20'd74, -20'd38, 20'd170, 20'd67, 20'd83, 20'd117, -20'd39, -20'd96, 20'd79, -20'd157, -20'd221, 20'd19, 20'd71, 20'd153, 20'd43, -20'd165, -20'd71, 20'd167, -20'd34, -20'd162, -20'd210, 20'd51};
