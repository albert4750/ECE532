localparam bit signed [0:146][7:0] Input6 = '{-112, -123, -88, 55, 29, 53, -106, -27, -105, 123, -6, 36, 107, 59, -94, 70, 6, -40, -52, -111, -33, -80, -91, -128, 74, -15, -20, -124, -33, 60, -1, -118, -99, -31, -23, 112, -115, -109, -87, 76, 44, -77, -21, 16, 120, 126, 114, 37, -114, 36, -14, 4, 114, -81, 0, -79, 37, 126, 75, -84, -59, -24, 110, -112, -112, -118, -123, 23, 47, -61, 38, 112, -110, -34, 80, -97, 42, -81, -107, 97, -73, -54, -20, -97, -45, -62, 19, 31, -14, -109, -89, 39, -67, -31, 44, 116, 108, 54, 94, -6, 103, 62, 76, 16, -48, 126, 6, 68, -83, 84, 122, 30, -52, -5, 53, 33, -38, 18, 6, -8, 2, 26, 110, -103, -115, 63, 91, -66, -71, -91, 45, 21, -21, 120, -59, 121, -79, -103, -116, -76, -58, 47, 125, -55, 10, -56, 90};
