localparam bit signed [0:2][47:0] Bias3 = '{48'd39088, -48'd90262, -48'd32497};
