localparam bit signed [0:7][47:0] Bias2 = '{48'd91918, -48'd146106, 48'd8658, 48'd180660, -48'd102780, -48'd121131, -48'd160817, -48'd51809};
