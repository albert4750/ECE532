localparam bit signed [0:7][47:0] Bias2 = '{48'd590311, 48'd591275, 48'd168954, 48'd433220, 48'd24212, 48'd425827, 48'd209602, 48'd433244};
