localparam bit signed [0:7][47:0] Bias1 = '{48'd4674, 48'd273918, -48'd29840, 48'd474992, -48'd108571, 48'd505490, 48'd749931, 48'd320401};
