localparam bit signed [0:15][7:0] Output4 = '{-34, 36, -12, 33, -48, -39, 41, -99, -124, 15, -76, -38, 91, -46, 68, -13};
