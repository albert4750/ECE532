localparam bit signed [0:7][47:0] Bias2 = '{48'd232707, -48'd242058, -48'd209802, 48'd227373, -48'd198352, 48'd95453, 48'd21432, 48'd203679};
