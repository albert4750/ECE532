localparam bit signed [0:63][0:2][0:8][0:8][24:0] Weight1 = '{
    '{'{'{-25'd193369, -25'd4756886, -25'd4447495, 25'd502760, -25'd2707171, 25'd2127063, -25'd696130, 25'd696130, -25'd3480648}, '{25'd502760, 25'd1044194, 25'd1701650, 25'd541434, -25'd3055235, -25'd2629823, -25'd3132583, 25'd3248605, 25'd2436454}, '{-25'd4795559, 25'd966847, -25'd386739, -25'd4331473, 25'd4602190, -25'd3480648, 25'd502760, 25'd2513801, -25'd1817672}, '{25'd1895019, -25'd1546955, 25'd3248605, 25'd4447495, -25'd425413, -25'd1198890, 25'd3132583, -25'd1662976, 25'd1430933}, '{-25'd1740324, -25'd1237564, -25'd4292799, 25'd464086, -25'd3944734, -25'd1198890, -25'd3441974, -25'd3287279, -25'd1121542}, '{25'd4640864, 25'd928173, 25'd4331473, 25'd1353585, 25'd2436454, 25'd3441974, -25'd232043, 25'd812151, -25'd4524842}, '{-25'd4640864, 25'd3867387, -25'd3325953, 25'd4138104, -25'd2629823, 25'd2629823, -25'd38674, -25'd4060756, 25'd77348}, '{25'd77348, -25'd2204410, 25'd2475127, -25'd4756886, 25'd3635343, -25'd2165737, 25'd2127063, 25'd1778998, 25'd3828713}, '{25'd1276238, 25'd3519322, -25'd502760, -25'd1585629, 25'd2707171, 25'd1392259, -25'd3016562, 25'd1701650, 25'd3093909}}, '{'{25'd2745845, -25'd4254125, -25'd773477, 25'd2784518, 25'd1972367, 25'd2127063, -25'd3287279, -25'd3209931, 25'd3790039}, '{-25'd928173, 25'd309391, 25'd2591149, 25'd1972367, -25'd541434, 25'd2861866, 25'd1895019, 25'd657456, -25'd1198890}, '{-25'd2939214, -25'd580108, -25'd4718212, -25'd812151, -25'd580108, 25'd3055235, -25'd348065, 25'd580108, 25'd2900540}, '{-25'd928173, 25'd2591149, -25'd4138104, -25'd2359106, -25'd3983408, -25'd4292799, -25'd1276238, 25'd2900540, -25'd3325953}, '{-25'd3055235, 25'd2977888, 25'd3519322, 25'd3325953, -25'd3248605, -25'd4138104, -25'd3596670, 25'd1740324, -25'd1353585}, '{-25'd3364626, 25'd348065, -25'd2900540, 25'd1624302, 25'd3364626, -25'd2591149, 25'd3209931, -25'd4911581, 25'd2049715}, '{25'd2281758, 25'd1160216, -25'd2397780, -25'd2745845, 25'd154695, 25'd154695, 25'd2475127, 25'd2243084, -25'd1585629}, '{25'd2823192, 25'd2552475, 25'd2668497, -25'd3983408, 25'd966847, 25'd270717, 25'd541434, 25'd1817672, 25'd309391}, '{25'd0, 25'd2397780, 25'd1701650, -25'd812151, -25'd3209931, 25'd38674, 25'd4331473, 25'd4718212, 25'd4254125}}, '{'{25'd4138104, -25'd2049715, 25'd3712691, 25'd928173, 25'd3751365, 25'd1314911, 25'd502760, -25'd3093909, -25'd4408821}, '{25'd348065, -25'd3790039, -25'd2900540, 25'd2165737, -25'd3906061, -25'd541434, 25'd928173, -25'd2397780, 25'd232043}, '{25'd3055235, -25'd1701650, -25'd734803, 25'd1237564, -25'd2243084, 25'd2977888, 25'd1469607, -25'd3674017, 25'd2397780}, '{25'd3557996, -25'd889499, 25'd1933693, -25'd2861866, 25'd2281758, 25'd4331473, -25'd4331473, -25'd541434, 25'd2977888}, '{-25'd3867387, 25'd1160216, -25'd4099430, -25'd1469607, -25'd4370147, -25'd3944734, 25'd2475127, -25'd4950255, -25'd3596670}, '{-25'd2127063, 25'd1082868, -25'd4447495, 25'd4679538, 25'd696130, 25'd2707171, -25'd4563516, -25'd348065, 25'd232043}, '{-25'd3055235, 25'd1082868, 25'd4060756, 25'd2977888, -25'd3132583, -25'd2900540, 25'd1121542, -25'd3364626, 25'd3055235}, '{-25'd2745845, -25'd3906061, 25'd4370147, -25'd2088389, -25'd1972367, -25'd270717, -25'd3983408, -25'd2243084, 25'd502760}, '{-25'd1701650, 25'd4022082, -25'd2707171, 25'd3751365, -25'd2436454, -25'd3751365, -25'd928173, -25'd3557996, 25'd3171257}}},
    '{'{'{-25'd2478249, 25'd3318333, -25'd294029, 25'd966097, -25'd4032404, 25'd4074409, 25'd2562257, -25'd546055, 25'd2856286}, '{-25'd672067, -25'd1512152, -25'd882088, 25'd4620463, 25'd1848185, 25'd4032404, -25'd3822383, 25'd2100211, -25'd504051}, '{-25'd3318333, 25'd4956497, -25'd1302131, -25'd3864388, 25'd4788480, 25'd4200421, -25'd2100211, 25'd4284430, -25'd3444345}, '{25'd3990400, -25'd3948396, -25'd3066307, 25'd2730274, 25'd2226223, -25'd1974198, 25'd1512152, -25'd84008, -25'd2688270}, '{25'd1932194, -25'd126013, 25'd4956497, 25'd5334535, -25'd3864388, 25'd3486350, -25'd2898291, -25'd2940295, -25'd2940295}, '{25'd3402341, 25'd2016202, 25'd1722173, 25'd3570358, 25'd798080, -25'd462046, 25'd5124514, 25'd5040505, -25'd924093}, '{-25'd1932194, 25'd1092110, -25'd4410442, 25'd2100211, 25'd3318333, -25'd630063, 25'd546055, 25'd2562257, 25'd1554156}, '{25'd3360337, -25'd2940295, 25'd504051, 25'd2478249, -25'd2562257, 25'd1386139, 25'd1764177, 25'd210021, -25'd1596160}, '{25'd504051, 25'd4704472, 25'd4914493, 25'd4200421, -25'd168017, 25'd168017, 25'd3402341, 25'd1806181, 25'd4074409}}, '{'{-25'd2478249, 25'd3360337, 25'd4536455, -25'd2982299, -25'd3570358, 25'd168017, -25'd3234324, 25'd4410442, -25'd3864388}, '{-25'd168017, 25'd2898291, -25'd4578459, -25'd3360337, 25'd2436244, -25'd588059, -25'd2772278, 25'd126013, 25'd798080}, '{-25'd4200421, -25'd2226223, 25'd2814282, 25'd3108312, -25'd3864388, 25'd756076, -25'd3738375, -25'd336034, -25'd2520253}, '{25'd2310232, -25'd882088, -25'd3906392, -25'd882088, -25'd1302131, 25'd1848185, 25'd1848185, 25'd3528354, -25'd966097}, '{25'd2982299, -25'd2184219, 25'd168017, -25'd2184219, -25'd588059, 25'd4830484, -25'd294029, 25'd4074409, -25'd3822383}, '{-25'd3738375, -25'd3150316, -25'd1974198, -25'd2814282, 25'd5082510, -25'd4662468, -25'd1302131, 25'd1092110, -25'd3402341}, '{25'd2982299, -25'd4872489, 25'd3024303, 25'd2184219, 25'd4536455, -25'd4788480, -25'd1050105, -25'd462046, 25'd1008101}, '{-25'd3822383, 25'd252025, 25'd2898291, -25'd3738375, 25'd4074409, 25'd4032404, -25'd3234324, 25'd1596160, -25'd1470147}, '{25'd3024303, 25'd462046, -25'd1806181, -25'd3192320, -25'd4536455, -25'd336034, -25'd1176118, 25'd4662468, -25'd1050105}}, '{'{25'd2268227, 25'd4914493, -25'd1470147, 25'd4830484, -25'd1722173, -25'd3486350, -25'd3234324, -25'd966097, 25'd2226223}, '{-25'd4326434, 25'd1932194, 25'd1134114, -25'd42004, 25'd42004, -25'd1596160, 25'd4242425, 25'd4116413, -25'd546055}, '{25'd2814282, -25'd1092110, -25'd1050105, 25'd798080, -25'd1806181, -25'd2772278, -25'd3948396, -25'd42004, 25'd2226223}, '{25'd2814282, -25'd504051, 25'd4704472, 25'd5166518, 25'd4746476, -25'd1932194, 25'd1848185, 25'd4410442, 25'd1806181}, '{25'd588059, 25'd2310232, 25'd1680168, 25'd5292531, 25'd4662468, 25'd1596160, 25'd2184219, -25'd3570358, -25'd798080}, '{25'd1512152, -25'd2268227, -25'd2520253, -25'd2058206, 25'd2394240, 25'd5208522, -25'd2562257, 25'd4494451, -25'd3654366}, '{25'd3360337, 25'd2436244, 25'd126013, -25'd2856286, -25'd588059, -25'd126013, 25'd2520253, 25'd4326434, 25'd1764177}, '{25'd378038, 25'd4872489, 25'd2142215, -25'd84008, 25'd1470147, -25'd252025, -25'd4620463, -25'd3444345, -25'd2058206}, '{25'd2226223, 25'd1050105, -25'd1554156, 25'd2436244, -25'd3234324, -25'd4368438, -25'd2478249, -25'd1512152, -25'd378038}}},
    '{'{'{25'd3147800, -25'd3893332, -25'd1573900, 25'd2526524, 25'd4887374, -25'd4017587, -25'd1822411, 25'd3354892, 25'd3189218}, '{25'd828368, 25'd3479147, 25'd4680282, -25'd1905247, -25'd994042, -25'd1159716, -25'd1822411, -25'd3727658, -25'd2899290}, '{25'd3396311, 25'd1698155, 25'd3313474, -25'd1739574, 25'd2733616, 25'd2526524, -25'd2278013, 25'd2319432, 25'd3520566}, '{25'd2236595, 25'd662695, 25'd3810495, -25'd4680282, -25'd2567942, -25'd911205, 25'd1408226, 25'd2816453, -25'd2278013}, '{-25'd3064963, 25'd2650779, -25'd745532, -25'd5094466, -25'd5011629, 25'd621276, -25'd704113, -25'd2816453, 25'd3479147}, '{25'd1159716, 25'd3354892, 25'd1863829, -25'd828368, -25'd4473190, 25'd538439, 25'd3064963, -25'd3479147, 25'd3023545}, '{-25'd3354892, 25'd3851913, -25'd4928792, 25'd2029503, -25'd124255, -25'd5094466, -25'd1325389, -25'd828368, 25'd1283971}, '{-25'd2692197, -25'd1366808, -25'd2236595, -25'd4017587, -25'd869787, 25'd2982126, 25'd4680282, 25'd2775034, -25'd372766}, '{25'd2195176, 25'd3810495, 25'd1201134, 25'd1573900, -25'd1573900, -25'd2029503, 25'd3147800, 25'd4183261, -25'd3437729}}, '{'{25'd4307516, 25'd1532482, 25'd4763119, 25'd2940708, -25'd1366808, 25'd331347, -25'd3686240, 25'd1988084, 25'd4348934}, '{-25'd1408226, 25'd414184, 25'd2360850, 25'd3520566, -25'd4183261, 25'd2485105, 25'd1905247, -25'd1532482, 25'd3769076}, '{25'd3893332, 25'd1118297, -25'd1366808, 25'd4100424, 25'd1822411, -25'd745532, -25'd1656737, 25'd3189218, 25'd2443687}, '{25'd3561984, -25'd2567942, 25'd1905247, 25'd2153758, 25'd3189218, -25'd2195176, -25'd5094466, -25'd1076879, -25'd786950}, '{-25'd3603403, -25'd1739574, -25'd3603403, -25'd1325389, -25'd3230637, -25'd2278013, 25'd2940708, 25'd2567942, -25'd1491063}, '{-25'd3396311, -25'd3230637, 25'd1739574, 25'd2650779, -25'd1822411, -25'd5135884, 25'd3479147, -25'd1159716, -25'd2899290}, '{-25'd1159716, 25'd2360850, 25'd124255, 25'd2982126, -25'd5218721, 25'd3851913, 25'd1573900, 25'd455603, -25'd4141842}, '{-25'd2153758, 25'd3147800, 25'd455603, -25'd3851913, 25'd3934750, -25'd2195176, -25'd3851913, 25'd2195176, -25'd4307516}, '{25'd3479147, -25'd372766, 25'd1905247, 25'd1076879, 25'd786950, 25'd3934750, -25'd4845955, 25'd3561984, -25'd4348934}}, '{'{-25'd4431771, -25'd1491063, -25'd704113, 25'd869787, -25'd786950, 25'd41418, 25'd2733616, -25'd1573900, -25'd1283971}, '{25'd4017587, 25'd2692197, -25'd538439, 25'd2650779, 25'd3023545, 25'd289929, 25'd3603403, -25'd4638863, -25'd2816453}, '{-25'd828368, 25'd1863829, -25'd3561984, 25'd3851913, -25'd828368, -25'd1325389, 25'd2485105, -25'd165674, -25'd1449645}, '{-25'd248511, -25'd2567942, 25'd621276, -25'd5011629, 25'd2526524, -25'd911205, 25'd2567942, -25'd1408226, -25'd3893332}, '{-25'd455603, 25'd4431771, -25'd662695, -25'd124255, 25'd3520566, -25'd828368, 25'd2733616, 25'd4059005, -25'd1573900}, '{25'd1946666, -25'd3354892, 25'd4307516, 25'd3396311, -25'd207092, -25'd579858, -25'd3189218, -25'd2153758, 25'd2733616}, '{25'd3644821, 25'd3106382, -25'd4680282, -25'd4307516, -25'd5301558, -25'd2692197, 25'd3023545, -25'd3313474, -25'd3727658}, '{-25'd2319432, 25'd4473190, 25'd1573900, 25'd2402268, 25'd1656737, 25'd331347, 25'd3354892, 25'd1242553, 25'd3644821}, '{-25'd4970211, -25'd3934750, 25'd3064963, -25'd2775034, 25'd704113, -25'd1325389, -25'd3272055, -25'd3769076, -25'd2692197}}},
    '{'{'{-25'd912378, 25'd608252, -25'd3779850, -25'd1998542, 25'd4909461, -25'd260679, 25'd4822568, 25'd912378, -25'd3041259}, '{-25'd4779121, 25'd2650240, -25'd3910190, 25'd738591, -25'd1303397, -25'd4648781, -25'd3997083, -25'd4952907, 25'd217233}, '{-25'd1390290, 25'd2476454, 25'd260679, -25'd2997812, -25'd2215774, 25'd4127423, -25'd4909461, -25'd3823297, 25'd3606064}, '{-25'd2259221, -25'd173786, 25'd2606793, -25'd2997812, 25'd2563347, 25'd4040530, 25'd4170869, 25'd3432278, 25'd1129610}, '{25'd4561888, -25'd3953636, -25'd4388102, -25'd4605335, 25'd4344655, -25'd1955095, 25'd1086164, 25'd4561888, -25'd3475724}, '{25'd1564076, -25'd1129610, -25'd4127423, 25'd4431549, -25'd260679, -25'd608252, -25'd1955095, 25'd4474995, 25'd3953636}, '{-25'd86893, 25'd521359, -25'd304126, 25'd2259221, -25'd1173057, -25'd3388831, -25'd2824026, 25'd4561888, 25'd1607523}, '{-25'd1737862, 25'd1173057, -25'd3866743, -25'd2476454, 25'd3910190, 25'd4040530, -25'd1390290, -25'd3692957, -25'd521359}, '{-25'd4822568, -25'd4127423, 25'd130340, 25'd217233, -25'd3258492, 25'd4518442, 25'd260679, -25'd2997812, 25'd1607523}}, '{'{-25'd3779850, 25'd2867473, -25'd955824, 25'd2910919, -25'd2476454, 25'd3475724, -25'd2476454, -25'd1824755, -25'd5474266}, '{-25'd2650240, -25'd1216504, 25'd3171598, -25'd2737133, 25'd2910919, 25'd782038, 25'd1694416, -25'd4735674, -25'd1390290}, '{25'd3823297, 25'd1998542, 25'd1955095, -25'd3606064, -25'd2954366, -25'd3953636, -25'd5517712, -25'd5561159, -25'd912378}, '{25'd3823297, 25'd1824755, -25'd955824, -25'd5430819, 25'd1520629, 25'd3997083, 25'd2997812, -25'd5126693, 25'd391019}, '{25'd4214316, 25'd2824026, 25'd2259221, 25'd1129610, 25'd4127423, 25'd2824026, -25'd1477183, 25'd260679, 25'd1737862}, '{-25'd3128152, 25'd2433007, 25'd3823297, -25'd4214316, 25'd521359, -25'd1911648, 25'd1390290, 25'd2433007, 25'd1129610}, '{25'd2476454, -25'd2389561, -25'd3606064, -25'd2780579, -25'd3171598, -25'd955824, 25'd477912, 25'd3475724, -25'd2910919}, '{-25'd4127423, -25'd4909461, -25'd1042717, -25'd1998542, 25'd2867473, 25'd3388831, -25'd347572, -25'd3779850, 25'd4301209}, '{-25'd4214316, 25'd1911648, 25'd347572, 25'd2346114, -25'd2302667, 25'd782038, -25'd86893, 25'd2476454, 25'd3562617}}, '{'{25'd868931, -25'd1477183, -25'd1694416, -25'd4561888, -25'd3736404, -25'd4692228, -25'd1390290, -25'd2563347, 25'd3736404}, '{-25'd1433736, -25'd695145, -25'd4214316, -25'd5474266, 25'd2476454, 25'd1433736, -25'd4648781, 25'd4040530, 25'd2519900}, '{25'd1607523, 25'd868931, -25'd5300480, -25'd5561159, 25'd477912, -25'd1520629, 25'd564805, -25'd3866743, 25'd651698}, '{25'd1216504, -25'd2606793, -25'd651698, 25'd2476454, -25'd173786, -25'd4692228, -25'd3041259, -25'd3171598, 25'd3779850}, '{25'd1259950, -25'd4779121, -25'd3866743, 25'd2824026, -25'd4474995, 25'd1346843, 25'd4474995, -25'd2606793, 25'd3128152}, '{-25'd2650240, -25'd2259221, 25'd2346114, 25'd4170869, 25'd1216504, 25'd3866743, 25'd1433736, 25'd4301209, 25'd2041988}, '{-25'd130340, -25'd2693686, -25'd3432278, 25'd1303397, 25'd651698, -25'd1216504, -25'd1998542, -25'd3562617, -25'd3345385}, '{-25'd3258492, 25'd695145, 25'd43447, 25'd3301938, -25'd3866743, 25'd4083976, -25'd391019, -25'd1824755, -25'd1781309}, '{25'd1390290, -25'd5126693, -25'd2389561, -25'd86893, -25'd868931, -25'd825485, 25'd2867473, 25'd1259950, -25'd825485}}},
    '{'{'{-25'd1491475, 25'd3728686, -25'd2747453, 25'd3296944, -25'd2629705, 25'd4749169, -25'd3218445, 25'd2472708, 25'd3964182}, '{-25'd2708204, -25'd1883968, 25'd1923217, 25'd627989, -25'd4395925, -25'd1491475, 25'd902735, -25'd1373727, -25'd5023914}, '{-25'd4317426, -25'd1020483, 25'd2825952, -25'd1412976, 25'd745737, -25'd4160429, 25'd3610938, 25'd1962466, 25'd2119464}, '{-25'd2354960, -25'd2433458, 25'd1412976, 25'd1295228, 25'd2708204, -25'd2786702, 25'd1059732, 25'd784987, 25'd1020483}, '{-25'd1177480, 25'd4945416, 25'd4474424, 25'd1216729, -25'd470992, 25'd2001716, 25'd2276461, 25'd1923217, -25'd2080214}, '{25'd1138231, 25'd3689437, -25'd4042681, 25'd784987, 25'd1844719, -25'd588740, -25'd2040965, 25'd392493, -25'd2276461}, '{-25'd4788418, 25'd706488, -25'd4081930, 25'd2982949, -25'd2119464, -25'd902735, -25'd4592172, -25'd2865201, -25'd392493}, '{25'd1569973, 25'd588740, -25'd2786702, -25'd2904450, 25'd3924933, -25'd2433458, -25'd510241, -25'd4238928, -25'd3022198}, '{-25'd1491475, 25'd2629705, 25'd824236, 25'd3179196, -25'd1138231, 25'd3414692, -25'd981233, 25'd4709920, 25'd4356676}}, '{'{25'd1805469, 25'd4395925, 25'd4356676, 25'd3218445, 25'd2825952, 25'd941984, 25'd2865201, -25'd2040965, 25'd3414692}, '{25'd2315710, 25'd549491, -25'd1098981, -25'd627989, -25'd2433458, -25'd2747453, 25'd1412976, 25'd39249, -25'd824236}, '{-25'd2511957, 25'd3022198, 25'd1177480, 25'd1569973, -25'd2080214, 25'd470992, -25'd2825952, 25'd2040965, 25'd1059732}, '{-25'd3885684, 25'd1138231, 25'd549491, 25'd1609223, 25'd2747453, 25'd1177480, 25'd510241, -25'd1138231, -25'd1844719}, '{25'd353244, -25'd1648472, -25'd745737, 25'd235496, 25'd392493, -25'd1766220, 25'd4199678, 25'd4866917, 25'd4199678}, '{-25'd4631421, -25'd3924933, -25'd4042681, 25'd1216729, 25'd2629705, -25'd1452225, 25'd3061448, 25'd706488, 25'd1923217}, '{25'd470992, -25'd4788418, 25'd0, -25'd470992, 25'd2786702, 25'd4631421, 25'd2315710, 25'd1805469, 25'd1569973}, '{-25'd4709920, 25'd3296944, -25'd4081930, 25'd1805469, 25'd2825952, -25'd353244, 25'd1805469, -25'd4513673, -25'd3610938}, '{-25'd3767936, 25'd2943700, 25'd4356676, -25'd1530724, -25'd4670670, 25'd1020483, -25'd4631421, 25'd2237212, 25'd863485}}, '{'{-25'd39249, -25'd3571689, -25'd4081930, 25'd1726971, -25'd2394209, 25'd3610938, 25'd2511957, -25'd4945416, 25'd2354960}, '{25'd2943700, -25'd3924933, -25'd1962466, 25'd2708204, 25'd4199678, -25'd1491475, 25'd4238928, 25'd510241, -25'd4395925}, '{25'd4552922, 25'd274745, -25'd4121180, -25'd549491, -25'd549491, 25'd1844719, -25'd2354960, 25'd1962466, -25'd4709920}, '{25'd2119464, -25'd1059732, 25'd2904450, -25'd1766220, -25'd235496, 25'd3453941, 25'd4552922, -25'd2158713, 25'd2982949}, '{-25'd3650188, 25'd4042681, -25'd3885684, -25'd4317426, -25'd3767936, 25'd235496, 25'd4513673, 25'd981233, 25'd1962466}, '{-25'd2982949, 25'd1098981, 25'd3257694, 25'd2315710, -25'd274745, -25'd1530724, 25'd4356676, 25'd1216729, 25'd2394209}, '{-25'd3807185, 25'd4199678, -25'd4866917, 25'd470992, -25'd3728686, 25'd4709920, -25'd1177480, -25'd2354960, -25'd4906166}, '{-25'd941984, 25'd274745, -25'd353244, 25'd3139946, -25'd941984, 25'd1569973, -25'd549491, -25'd2237212, 25'd2040965}, '{-25'd1098981, -25'd2080214, -25'd3571689, 25'd3375442, 25'd4199678, -25'd274745, -25'd2511957, 25'd2904450, 25'd2668954}}},
    '{'{'{-25'd1932948, -25'd3084492, -25'd4400541, 25'd2056328, 25'd3619137, -25'd2426467, -25'd1727315, 25'd329012, 25'd4153782}, '{-25'd2426467, 25'd4729554, 25'd4318288, 25'd4194909, 25'd4647301, -25'd1809568, -25'd3742516, 25'd3536884, 25'd123380}, '{-25'd2919985, -25'd1562809, 25'd4112655, 25'd411266, -25'd123380, 25'd5140819, -25'd2590973, -25'd2878859, 25'd3660263}, '{-25'd2467593, -25'd4194909, -25'd82253, -25'd1932948, 25'd4441668, 25'd3865896, -25'd82253, 25'd1233797, -25'd534645}, '{25'd3248998, 25'd1192670, -25'd2056328, 25'd3166745, 25'd2590973, 25'd2426467, -25'd534645, 25'd1357176, -25'd4523921}, '{-25'd2220834, 25'd4770680, 25'd4236035, 25'd2138581, 25'd616898, -25'd2961112, 25'd82253, -25'd2549846, -25'd1645062}, '{25'd3166745, 25'd2426467, 25'd4688427, 25'd987037, -25'd3331251, -25'd616898, -25'd1521682, 25'd4277162, -25'd1480556}, '{25'd1727315, -25'd1562809, 25'd3290124, -25'd4482794, 25'd699151, 25'd3948149, -25'd1028164, -25'd3701390, -25'd1521682}, '{25'd3331251, -25'd2878859, -25'd1233797, -25'd4811807, 25'd3989276, 25'd1069290, -25'd2385340, -25'd41127, -25'd3454631}}, '{'{25'd329012, 25'd2015201, 25'd4236035, 25'd2220834, -25'd4729554, 25'd2385340, 25'd1398303, -25'd1974075, -25'd4482794}, '{25'd2097454, 25'd4194909, 25'd3290124, 25'd5017440, 25'd1850695, 25'd3331251, -25'd658025, 25'd329012, -25'd1398303}, '{-25'd4112655, -25'd3290124, -25'd1274923, -25'd3454631, -25'd1974075, -25'd3207871, 25'd2344214, 25'd0, 25'd3536884}, '{25'd904784, -25'd2220834, 25'd3865896, -25'd1686189, 25'd1645062, -25'd1069290, -25'd1151544, 25'd2755479, -25'd987037}, '{25'd3454631, -25'd3413504, -25'd3372377, -25'd3413504, 25'd3536884, 25'd3166745, 25'd1768442, 25'd4729554, 25'd4359415}, '{25'd2919985, 25'd3660263, -25'd1069290, 25'd3454631, 25'd287886, 25'd1974075, -25'd3989276, -25'd4565047, -25'd4071529}, '{-25'd699151, 25'd1192670, 25'd3989276, -25'd1686189, 25'd2919985, 25'd1110417, -25'd3701390, 25'd4030402, -25'd534645}, '{-25'd2919985, -25'd3495757, -25'd2261960, -25'd4606174, 25'd1233797, -25'd740278, 25'd1316050, -25'd3372377, 25'd4400541}, '{25'd41127, 25'd1316050, 25'd411266, -25'd287886, -25'd3865896, -25'd287886, 25'd4441668, 25'd3619137, 25'd2179707}}, '{'{-25'd1316050, -25'd1316050, 25'd2919985, 25'd2261960, -25'd863658, -25'd904784, -25'd3454631, 25'd3331251, 25'd575772}, '{-25'd1562809, -25'd3002238, -25'd4688427, -25'd2878859, -25'd205633, 25'd2344214, 25'd3331251, -25'd1686189, -25'd1562809}, '{-25'd4194909, 25'd3783643, 25'd2755479, -25'd863658, 25'd2179707, 25'd863658, 25'd3948149, 25'd1809568, -25'd3495757}, '{-25'd2590973, -25'd4030402, 25'd3125618, 25'd4112655, 25'd5223072, 25'd5140819, 25'd3207871, -25'd1274923, 25'd987037}, '{-25'd1809568, -25'd2220834, -25'd1357176, 25'd1069290, 25'd5223072, 25'd3989276, 25'd1192670, -25'd3742516, 25'd2919985}, '{-25'd4647301, 25'd3290124, 25'd1645062, 25'd4194909, -25'd1028164, 25'd1768442, 25'd3824770, 25'd287886, 25'd4976313}, '{25'd4811807, 25'd1274923, 25'd3372377, 25'd3907023, 25'd1398303, 25'd2015201, -25'd4236035, -25'd452392, 25'd575772}, '{-25'd2344214, -25'd781405, -25'd699151, 25'd4194909, -25'd4606174, 25'd3865896, 25'd1603936, 25'd4441668, 25'd1110417}, '{25'd4194909, -25'd4729554, 25'd1974075, 25'd575772, 25'd1603936, 25'd2673226, 25'd2467593, -25'd4318288, 25'd2344214}}},
    '{'{'{25'd4223761, -25'd3620367, 25'd2852410, -25'd6527631, -25'd5046572, -25'd3016972, -25'd3126681, -25'd4662594, -25'd4662594}, '{25'd877665, 25'd5265988, 25'd3346097, -25'd4827156, 25'd1590767, -25'd3071826, -25'd219416, 25'd1865038, 25'd1426205}, '{25'd2084454, 25'd713103, -25'd5869383, -25'd1426205, -25'd1426205, -25'd4662594, -25'd164562, -25'd274270, -25'd2249016}, '{25'd932519, -25'd1590767, -25'd1810183, 25'd713103, -25'd4443178, -25'd987373, 25'd4498032, 25'd1042227, -25'd4443178}, '{-25'd1481059, -25'd4991718, -25'd1590767, -25'd4662594, -25'd383978, 25'd822811, 25'd4607740, -25'd3016972, 25'd1919892}, '{-25'd3784929, -25'd4991718, 25'd548540, -25'd3400951, 25'd1151935, -25'd767957, 25'd5156280, 25'd2523286, -25'd493686}, '{25'd383978, -25'd1535913, -25'd219416, 25'd2303870, 25'd383978, 25'd5704821, 25'd5265988, -25'd3236389, 25'd822811}, '{25'd4991718, -25'd164562, -25'd2084454, -25'd1426205, 25'd54854, -25'd2358724, -25'd2797556, -25'd3784929, -25'd877665}, '{25'd109708, -25'd3400951, 25'd5704821, 25'd2797556, 25'd4114053, -25'd1426205, -25'd5320842, -25'd1316497, -25'd987373}}, '{'{25'd4388324, -25'd2852410, -25'd2358724, -25'd4662594, 25'd329124, 25'd329124, 25'd1316497, 25'd383978, 25'd1042227}, '{25'd4443178, 25'd2084454, -25'd1919892, 25'd2797556, -25'd6198507, 25'd2907264, 25'd3675221, 25'd1535913, 25'd2962118}, '{25'd2084454, -25'd1097081, -25'd274270, -25'd7021318, 25'd2358724, -25'd2687848, 25'd1151935, 25'd3894637, -25'd3510659}, '{25'd2962118, -25'd4827156, 25'd329124, -25'd5540258, -25'd1645621, 25'd3620367, 25'd4114053, 25'd4004345, 25'd2852410}, '{-25'd2029600, -25'd5211134, -25'd6308215, 25'd2907264, 25'd1865038, 25'd1042227, 25'd4772302, 25'd3346097, -25'd2029600}, '{-25'd5704821, -25'd3346097, -25'd2303870, -25'd2303870, 25'd5595113, 25'd3839783, 25'd4388324, 25'd329124, 25'd2852410}, '{-25'd3675221, 25'd3784929, -25'd1590767, 25'd1371351, 25'd4717448, 25'd109708, 25'd2742702, 25'd274270, 25'd2523286}, '{25'd548540, 25'd1810183, 25'd4936864, 25'd5101426, 25'd3894637, 25'd1535913, 25'd2194162, 25'd3291243, -25'd383978}, '{25'd3949491, -25'd2797556, 25'd1700475, 25'd3400951, 25'd3181535, -25'd3510659, 25'd2303870, -25'd438832, 25'd987373}}, '{'{25'd5485404, 25'd54854, 25'd2742702, -25'd1481059, 25'd2632994, 25'd438832, 25'd713103, 25'd164562, 25'd3839783}, '{25'd5156280, -25'd1974746, 25'd3236389, 25'd2194162, -25'd1810183, 25'd1974746, -25'd767957, 25'd3839783, -25'd1700475}, '{25'd4936864, 25'd164562, -25'd4827156, -25'd1426205, -25'd877665, 25'd2249016, -25'd987373, -25'd383978, 25'd932519}, '{-25'd2358724, -25'd4059199, -25'd4278615, -25'd6033945, -25'd5430550, -25'd3071826, -25'd3510659, -25'd2413578, -25'd3565513}, '{-25'd1755329, 25'd1755329, 25'd3346097, -25'd5375696, 25'd3565513, -25'd1426205, -25'd3784929, -25'd2523286, -25'd4223761}, '{-25'd2852410, -25'd1042227, 25'd54854, 25'd3730075, 25'd1919892, 25'd1261643, 25'd2139308, 25'd164562, -25'd4552886}, '{-25'd2907264, -25'd1590767, 25'd2249016, 25'd3016972, 25'd5265988, 25'd493686, -25'd2687848, 25'd4223761, -25'd1316497}, '{25'd109708, 25'd4388324, 25'd1261643, 25'd5759675, -25'd603394, -25'd2907264, 25'd2962118, 25'd658249, -25'd383978}, '{-25'd3620367, 25'd4278615, 25'd5485404, -25'd4333469, -25'd1590767, 25'd109708, -25'd4991718, -25'd5924237, 25'd658249}}},
    '{'{'{-25'd2605885, -25'd2124799, 25'd3086972, -25'd2886519, -25'd2245071, -25'd3247334, 25'd3888783, -25'd1483350, 25'd481087}, '{-25'd1322988, -25'd2686066, 25'd4129326, 25'd2084708, -25'd2405433, -25'd1804075, 25'd2766248, 25'd3568058, -25'd2525704}, '{-25'd881992, -25'd3768511, 25'd1643712, 25'd4289688, 25'd2164889, 25'd4650503, 25'd2204980, 25'd4129326, -25'd2565795}, '{25'd3006791, -25'd1804075, -25'd641449, -25'd2645976, 25'd761720, -25'd481087, -25'd841901, -25'd3527968, 25'd1964437}, '{-25'd3327515, -25'd4610413, 25'd3407696, -25'd3487877, -25'd3568058, 25'd4009054, 25'd1403169, 25'd1763984, 25'd4249598}, '{25'd2084708, -25'd2766248, 25'd1242807, -25'd681539, -25'd3327515, 25'd1282897, 25'd4169417, -25'd1242807, 25'd3086972}, '{25'd2124799, 25'd641449, -25'd1844165, 25'd1002264, -25'd440996, 25'd1443260, -25'd1804075, 25'd1042354, 25'd3287425}, '{-25'd4049145, 25'd2806338, -25'd2485614, 25'd4610413, -25'd2565795, 25'd2405433, 25'd3327515, -25'd3688330, 25'd3527968}, '{25'd1523441, 25'd4209507, -25'd40091, -25'd601358, 25'd440996, 25'd481087, 25'd1884256, -25'd4450050, -25'd2084708}}, '{'{25'd4730684, 25'd3167153, 25'd160362, 25'd1563531, -25'd601358, 25'd3247334, -25'd440996, 25'd2846429, 25'd4850956}, '{25'd2846429, 25'd2405433, -25'd1603622, -25'd1483350, 25'd2806338, -25'd3287425, 25'd4730684, 25'd1723893, -25'd962173}, '{25'd2766248, 25'd4931137, 25'd3287425, 25'd1042354, 25'd2966700, -25'd3768511, 25'd4289688, -25'd3247334, 25'd2445523}, '{25'd4089236, -25'd3207244, -25'd2645976, -25'd1483350, -25'd4329779, 25'd3808602, -25'd4329779, 25'd1282897, 25'd3487877}, '{-25'd3247334, -25'd3888783, -25'd80181, 25'd2605885, 25'd120272, 25'd962173, 25'd3527968, 25'd320724, 25'd1322988}, '{-25'd2164889, -25'd681539, -25'd4409960, 25'd4049145, -25'd561268, 25'd240543, 25'd5091499, -25'd1844165, -25'd1082445}, '{25'd160362, -25'd1723893, -25'd3287425, 25'd2525704, -25'd2044618, -25'd561268, 25'd3808602, 25'd4850956, 25'd4610413}, '{-25'd1122535, 25'd360815, 25'd561268, 25'd4850956, 25'd2806338, 25'd4850956, 25'd1763984, -25'd2605885, -25'd3127062}, '{25'd320724, 25'd1964437, -25'd1483350, -25'd4089236, 25'd2806338, -25'd2645976, -25'd922083, 25'd561268, -25'd3046881}}, '{'{-25'd1122535, 25'd2164889, -25'd4209507, 25'd601358, -25'd3768511, 25'd3407696, -25'd1844165, 25'd1322988, 25'd2766248}, '{-25'd2686066, 25'd841901, 25'd521177, -25'd1322988, -25'd4129326, -25'd4169417, 25'd1523441, -25'd1282897, 25'd0}, '{-25'd40091, 25'd4409960, 25'd400905, 25'd80181, 25'd4490141, -25'd280634, 25'd1964437, 25'd4730684, -25'd3086972}, '{25'd4450050, 25'd721630, -25'd400905, 25'd4490141, -25'd1964437, -25'd360815, -25'd1082445, -25'd4169417, -25'd3447787}, '{-25'd1804075, 25'd1322988, -25'd2084708, 25'd2886519, 25'd4209507, -25'd280634, 25'd1162626, 25'd3688330, 25'd1844165}, '{25'd1643712, -25'd3407696, -25'd3688330, -25'd2285161, 25'd3247334, 25'd721630, -25'd2365342, -25'd2445523, 25'd922083}, '{25'd2645976, -25'd721630, 25'd40091, 25'd3247334, -25'd3768511, -25'd4650503, -25'd801811, 25'd4730684, -25'd3207244}, '{25'd4409960, -25'd641449, -25'd1964437, -25'd3568058, -25'd1403169, -25'd4610413, 25'd3568058, -25'd3848692, -25'd440996}, '{-25'd3247334, -25'd962173, -25'd1162626, -25'd40091, 25'd4089236, 25'd2204980, -25'd2485614, 25'd2926610, 25'd2445523}}},
    '{'{'{25'd525557, -25'd565984, 25'd2263937, 25'd4770439, -25'd3840608, -25'd161710, 25'd1819235, -25'd1576670, -25'd3395906}, '{-25'd1091541, -25'd3598043, 25'd2021372, -25'd1293678, 25'd4608729, 25'd727694, -25'd808549, 25'd3598043, -25'd1495816}, '{-25'd404274, 25'd3678898, -25'd3032059, -25'd1334106, 25'd5134286, 25'd4568302, 25'd646839, -25'd1536243, -25'd2142655}, '{-25'd3072486, -25'd1980945, 25'd1455388, 25'd2061800, 25'd4244882, 25'd2263937, 25'd3193768, -25'd40427, -25'd1293678}, '{25'd2183082, 25'd1455388, 25'd0, -25'd3355478, -25'd4204455, 25'd4244882, -25'd485129, 25'd4891721, 25'd1657525}, '{25'd3759753, 25'd80855, 25'd80855, 25'd2829921, -25'd1495816, -25'd121282, 25'd2668212, 25'd0, 25'd727694}, '{25'd1131969, 25'd121282, -25'd2951204, 25'd4810866, 25'd4891721, -25'd2910776, -25'd2668212, -25'd970259, -25'd3193768}, '{-25'd1617098, -25'd1051114, -25'd1212823, -25'd1172396, 25'd5134286, -25'd646839, 25'd2183082, 25'd4608729, -25'd1940517}, '{25'd4810866, 25'd2263937, 25'd80855, -25'd3234196, 25'd687267, -25'd1617098, 25'd3759753, -25'd4285309, 25'd2344792}}, '{'{-25'd4487447, -25'd1697953, 25'd4285309, -25'd121282, 25'd2183082, -25'd1374533, 25'd1374533, 25'd4527874, -25'd2951204}, '{-25'd40427, -25'd161710, -25'd3395906, 25'd1212823, 25'd1940517, -25'd1212823, -25'd3476761, 25'd3759753, -25'd1212823}, '{25'd3759753, -25'd3840608, -25'd3234196, -25'd1778808, 25'd444702, -25'd40427, -25'd4487447, -25'd3638470, -25'd323420}, '{-25'd202137, 25'd2708639, 25'd2749066, 25'd5093858, -25'd1859663, 25'd808549, 25'd3193768, 25'd4689584, 25'd646839}, '{25'd2708639, -25'd2627784, -25'd4002317, 25'd4689584, 25'd2870349, 25'd848976, -25'd4325737, 25'd3678898, 25'd4244882}, '{25'd848976, 25'd1010686, -25'd40427, 25'd4285309, 25'd4972576, 25'd121282, 25'd848976, -25'd3759753, -25'd2466074}, '{25'd2466074, 25'd2021372, -25'd525557, 25'd646839, -25'd4002317, -25'd1738380, -25'd768122, 25'd1212823, -25'd1738380}, '{25'd3112913, -25'd4689584, -25'd4730011, -25'd1657525, 25'd3153341, 25'd1455388, 25'd4285309, -25'd282992, 25'd4891721}, '{-25'd1617098, 25'd3961890, -25'd4002317, 25'd2991631, -25'd3072486, -25'd3961890, 25'd0, 25'd2910776, 25'd3678898}}, '{'{25'd929831, 25'd3436333, 25'd525557, -25'd3112913, -25'd2546929, -25'd3274623, -25'd3193768, 25'd3395906, -25'd646839}, '{-25'd3234196, 25'd3274623, -25'd4042745, 25'd2789494, 25'd1819235, -25'd4204455, 25'd4608729, 25'd2991631, -25'd2385219}, '{25'd4042745, -25'd2385219, -25'd2870349, 25'd2627784, 25'd2021372, -25'd2991631, 25'd2991631, 25'd808549, -25'd2183082}, '{25'd4204455, 25'd3800180, -25'd4002317, -25'd768122, 25'd2627784, 25'd4447019, -25'd3153341, 25'd4932149, 25'd3800180}, '{-25'd242565, 25'd4325737, 25'd1091541, 25'd5093858, -25'd2102227, 25'd4972576, -25'd1334106, -25'd121282, 25'd1657525}, '{-25'd808549, -25'd1334106, -25'd2304365, -25'd1576670, -25'd161710, 25'd4608729, -25'd2385219, -25'd2102227, -25'd1253251}, '{-25'd1859663, -25'd2910776, 25'd727694, 25'd2910776, -25'd3598043, 25'd3598043, 25'd40427, -25'd4123600, 25'd161710}, '{25'd1617098, -25'd2587357, -25'd2304365, -25'd4568302, 25'd4002317, 25'd40427, 25'd3759753, 25'd525557, 25'd4527874}, '{-25'd2749066, 25'd1334106, -25'd3800180, 25'd1212823, 25'd4447019, 25'd3315051, -25'd2546929, -25'd4002317, 25'd1293678}}},
    '{'{'{25'd963066, -25'd4614690, 25'd521661, 25'd0, -25'd3049708, 25'd3170092, -25'd321022, 25'd3290475, 25'd1845876}, '{-25'd1564982, 25'd3852263, -25'd882810, -25'd1645237, 25'd2608303, -25'd2367537, 25'd2969453, -25'd1845876, 25'd4454179}, '{-25'd160511, -25'd200639, -25'd2688559, 25'd80255, 25'd2247154, -25'd3531241, -25'd240766, -25'd3731880, 25'd1805748}, '{25'd2608303, -25'd4654818, 25'd1003194, 25'd3892391, 25'd1645237, 25'd4614690, -25'd4213413, -25'd2768814, -25'd521661}, '{25'd1605110, 25'd2207026, 25'd4494307, 25'd3731880, 25'd3250347, -25'd120383, -25'd2608303, -25'd2247154, 25'd1966259}, '{25'd2046515, 25'd2487920, -25'd1364343, -25'd1444599, -25'd2327409, -25'd4173285, 25'd4052902, 25'd3049708, 25'd2969453}, '{-25'd3731880, -25'd1524854, 25'd280894, 25'd2247154, 25'd722299, -25'd882810, -25'd3731880, 25'd3932519, 25'd40128}, '{25'd3651625, -25'd280894, -25'd3812136, 25'd1805748, -25'd2126770, 25'd963066, -25'd3571369, -25'd4253541, 25'd3972647}, '{25'd1043321, 25'd240766, -25'd1564982, 25'd2166898, -25'd682172, 25'd682172, -25'd481533, -25'd1003194, 25'd3450986}}, '{'{-25'd1524854, 25'd2247154, -25'd120383, -25'd3531241, 25'd2648431, 25'd3852263, -25'd2487920, -25'd922938, 25'd3812136}, '{25'd1805748, -25'd3210219, -25'd3410858, 25'd0, 25'd0, 25'd4454179, 25'd1243960, 25'd3932519, -25'd3571369}, '{-25'd2929325, 25'd4614690, -25'd240766, 25'd3450986, -25'd2447792, -25'd3009581, -25'd3410858, 25'd2166898, 25'd4133157}, '{25'd3812136, -25'd3691752, 25'd4133157, -25'd4454179, -25'd1003194, 25'd1043321, -25'd80255, -25'd1805748, -25'd3129964}, '{-25'd3210219, 25'd4614690, 25'd1765621, 25'd1444599, -25'd842683, -25'd2969453, -25'd2126770, -25'd1243960, 25'd1524854}, '{25'd4253541, 25'd1484726, -25'd4454179, -25'd3290475, -25'd762427, -25'd3571369, -25'd561788, 25'd2046515, -25'd1926132}, '{-25'd3611497, 25'd682172, -25'd2768814, 25'd1605110, 25'd4454179, -25'd2046515, -25'd4775201, 25'd1364343, 25'd3651625}, '{-25'd2568176, 25'd3089836, -25'd2528048, 25'd682172, -25'd2046515, -25'd361150, -25'd4012774, -25'd802555, -25'd4012774}, '{-25'd4574563, 25'd682172, -25'd1444599, -25'd481533, -25'd3370730, 25'd3531241, 25'd120383, -25'd722299, 25'd642044}}, '{'{-25'd2166898, -25'd321022, -25'd3210219, -25'd401277, -25'd4654818, -25'd762427, 25'd521661, -25'd2046515, 25'd2608303}, '{25'd4213413, 25'd2969453, 25'd601916, -25'd40128, 25'd842683, -25'd2648431, -25'd3450986, -25'd2528048, 25'd3450986}, '{25'd3812136, -25'd922938, -25'd401277, -25'd2086643, -25'd1123577, -25'd2287281, 25'd722299, 25'd1805748, 25'd2648431}, '{25'd722299, -25'd4815329, -25'd5096223, 25'd1284088, -25'd2126770, 25'd2327409, -25'd4534435, 25'd2969453, 25'd361150}, '{-25'd2808942, -25'd2287281, -25'd2969453, -25'd4253541, 25'd1364343, 25'd3290475, 25'd642044, 25'd4414052, -25'd642044}, '{25'd1123577, 25'd762427, 25'd3089836, 25'd1765621, 25'd922938, -25'd2728686, -25'd3410858, 25'd1605110, -25'd963066}, '{25'd441405, -25'd4574563, -25'd4614690, 25'd3330603, -25'd1364343, -25'd1243960, -25'd240766, 25'd4654818, 25'd1564982}, '{-25'd2728686, -25'd882810, -25'd682172, 25'd4534435, -25'd4534435, -25'd4133157, -25'd1484726, -25'd4093030, 25'd601916}, '{-25'd722299, 25'd2969453, -25'd3691752, -25'd642044, 25'd2849070, -25'd3531241, -25'd1444599, 25'd2447792, 25'd3009581}}},
    '{'{'{-25'd2978254, -25'd386786, -25'd3481076, 25'd1972610, -25'd2823539, -25'd4796149, -25'd3016932, -25'd2668825, 25'd1585823}, '{-25'd4254648, -25'd2591467, -25'd2204681, 25'd4680113, 25'd773572, 25'd4486720, -25'd3442397, 25'd425465, 25'd3558433}, '{-25'd2127324, -25'd4796149, -25'd4873506, -25'd3713147, -25'd2784861, -25'd232072, -25'd2746182, 25'd3635790, 25'd3790505}, '{-25'd3481076, -25'd2552789, -25'd3983898, 25'd2978254, 25'd696215, -25'd386786, -25'd734894, 25'd580179, 25'd1972610}, '{-25'd3326361, 25'd3442397, -25'd4486720, 25'd1431109, -25'd3519754, 25'd966965, -25'd1469788, 25'd2978254, 25'd4641434}, '{-25'd2978254, 25'd3055611, 25'd4332005, 25'd3094290, 25'd2282039, -25'd1392430, -25'd1585823, 25'd2282039, 25'd1779216}, '{-25'd4448041, 25'd2088645, -25'd154714, -25'd1315073, -25'd2784861, 25'd1353752, -25'd3249004, -25'd1392430, -25'd77357}, '{25'd4641434, -25'd4950863, -25'd1044323, -25'd2243360, -25'd116036, -25'd3635790, -25'd4564077, -25'd4486720, 25'd38679}, '{-25'd4448041, 25'd1508466, -25'd1315073, 25'd3055611, -25'd502822, 25'd812251, 25'd2127324, -25'd4718792, 25'd3635790}}, '{'{25'd4448041, 25'd4564077, 25'd4641434, -25'd4680113, -25'd2552789, 25'd464143, -25'd4409363, 25'd348108, -25'd734894}, '{-25'd2707503, -25'd4718792, -25'd3171647, -25'd3132968, -25'd309429, -25'd812251, -25'd1624502, -25'd773572, 25'd2591467}, '{25'd1469788, -25'd1199037, -25'd270750, -25'd1199037, 25'd2978254, 25'd2668825, -25'd1779216, 25'd38679, -25'd3558433}, '{25'd1663181, -25'd2978254, -25'd1353752, -25'd3829183, -25'd2591467, -25'd3713147, 25'd386786, 25'd2746182, -25'd2823539}, '{25'd2746182, -25'd502822, -25'd541501, -25'd4834827, -25'd1856574, 25'd2630146, 25'd3790505, 25'd348108, 25'd1237716}, '{-25'd657537, 25'd1469788, 25'd2939575, 25'd3829183, 25'd889608, 25'd4138612, -25'd2127324, 25'd1431109, 25'd3016932}, '{25'd2784861, 25'd2088645, 25'd812251, -25'd2514110, -25'd1817895, 25'd2127324, 25'd77357, 25'd2668825, -25'd2243360}, '{-25'd3558433, 25'd2243360, 25'd1547145, 25'd1972610, -25'd2049967, -25'd1392430, -25'd3519754, 25'd2475432, -25'd4138612}, '{-25'd4641434, -25'd1508466, -25'd4680113, -25'd3558433, 25'd2668825, -25'd425465, -25'd2320717, -25'd2243360, 25'd734894}}, '{'{-25'd889608, 25'd850930, 25'd3519754, -25'd4796149, -25'd3790505, -25'd3867862, -25'd4641434, -25'd4409363, 25'd966965}, '{-25'd773572, 25'd1083001, -25'd464143, -25'd1972610, 25'd425465, 25'd1237716, 25'd116036, -25'd3983898, -25'd773572}, '{25'd1469788, 25'd2978254, 25'd4409363, 25'd3519754, 25'd4099934, -25'd3055611, 25'd1701859, 25'd386786, 25'd1817895}, '{25'd1392430, 25'd3094290, -25'd270750, 25'd2049967, -25'd1005644, 25'd3171647, -25'd3829183, -25'd4448041, -25'd734894}, '{-25'd3674469, 25'd1276394, 25'd3597112, 25'd3287683, -25'd812251, -25'd2011288, 25'd1431109, -25'd3558433, -25'd4718792}, '{-25'd1276394, 25'd4718792, -25'd3326361, -25'd3558433, -25'd2668825, -25'd1315073, -25'd2088645, -25'd4796149, 25'd3945219}, '{-25'd3635790, 25'd38679, 25'd1431109, -25'd4254648, 25'd3945219, 25'd1779216, -25'd2707503, 25'd3519754, 25'd3365040}, '{-25'd3635790, -25'd3132968, 25'd3829183, -25'd889608, -25'd734894, -25'd4293327, -25'd2978254, 25'd2591467, -25'd3326361}, '{-25'd2475432, -25'd2939575, 25'd2320717, 25'd4099934, -25'd2204681, -25'd502822, -25'd2320717, 25'd3867862, -25'd3210325}}},
    '{'{'{25'd3773835, -25'd3732364, -25'd580590, -25'd1866182, -25'd165883, 25'd3856776, 25'd1534416, 25'd4271483, -25'd373236}, '{25'd4810603, -25'd331766, 25'd3690893, 25'd705002, -25'd1410004, -25'd3442069, -25'd207354, 25'd0, -25'd3566481}, '{-25'd787944, 25'd3400598, 25'd4520308, 25'd2944421, -25'd3649423, 25'd1492946, -25'd3234716, 25'd4064130, -25'd82941}, '{25'd2654126, 25'd2363831, -25'd2032065, 25'd1949124, 25'd2529713, 25'd3566481, -25'd705002, 25'd1575887, -25'd2695596}, '{25'd2944421, -25'd1907653, 25'd995297, -25'd2778538, -25'd2197948, -25'd41471, 25'd373236, 25'd2778538, 25'd3400598}, '{25'd2280889, 25'd2571184, 25'd663531, 25'd2985891, -25'd207354, -25'd1327063, 25'd3317657, 25'd4976486, -25'd1119709}, '{25'd1575887, 25'd3981188, 25'd622061, -25'd456178, -25'd912356, -25'd4395896, 25'd1119709, 25'd4105601, 25'd4520308}, '{25'd4022659, 25'd4147071, 25'd2488243, 25'd2944421, 25'd3359128, 25'd2280889, -25'd456178, 25'd124412, -25'd290295}, '{-25'd2488243, -25'd3151774, 25'd1036768, 25'd3234716, 25'd1327063, -25'd2073536, 25'd3317657, -25'd2115006, 25'd4810603}}, '{'{25'd2239418, -25'd414707, 25'd3939718, -25'd2695596, -25'd2944421, 25'd165883, -25'd2073536, -25'd207354, -25'd1410004}, '{25'd1700299, 25'd1078239, 25'd539119, 25'd2363831, -25'd539119, 25'd2156477, 25'd1161180, -25'd1244121, -25'd1907653}, '{25'd1327063, 25'd4852073, 25'd1036768, -25'd1410004, -25'd1617358, 25'd3815306, 25'd2695596, -25'd3483540, 25'd1907653}, '{25'd1824711, 25'd3442069, 25'd290295, -25'd2944421, -25'd3981188, 25'd3110303, -25'd1617358, -25'd1410004, -25'd1244121}, '{-25'd4230013, 25'd1824711, -25'd1700299, -25'd3690893, 25'd995297, 25'd41471, 25'd4727661, 25'd1451475, -25'd4520308}, '{25'd663531, 25'd165883, -25'd787944, -25'd3773835, -25'd2032065, -25'd2322360, -25'd3276186, -25'd497649, 25'd1658829}, '{-25'd787944, -25'd373236, 25'd4976486, -25'd4520308, 25'd2820008, -25'd1410004, 25'd1368534, -25'd1451475, -25'd2529713}, '{25'd4644720, -25'd414707, 25'd746473, 25'd4354425, 25'd1119709, 25'd5142368, 25'd4810603, -25'd2446772, 25'd3981188}, '{25'd2902950, -25'd3981188, 25'd3483540, 25'd1617358, 25'd3525011, -25'd2695596, 25'd2944421, -25'd4312954, 25'd2239418}}, '{'{-25'd3690893, 25'd82941, 25'd1078239, -25'd2073536, -25'd2861479, -25'd2156477, 25'd124412, -25'd3317657, -25'd1824711}, '{-25'd4271483, 25'd663531, -25'd2032065, 25'd2197948, -25'd3317657, 25'd4852073, -25'd456178, -25'd3317657, -25'd3856776}, '{25'd953826, -25'd2197948, 25'd5059427, 25'd331766, 25'd4727661, -25'd2654126, 25'd4561778, -25'd2529713, -25'd1492946}, '{25'd290295, -25'd3773835, 25'd3193245, 25'd3815306, 25'd5266781, 25'd622061, 25'd2902950, 25'd2405301, 25'd4852073}, '{-25'd787944, 25'd1036768, -25'd2197948, -25'd3566481, 25'd1202651, 25'd5266781, 25'd5266781, 25'd3939718, 25'd3649423}, '{-25'd829414, -25'd4064130, 25'd2156477, 25'd4147071, -25'd2073536, 25'd3939718, -25'd2446772, 25'd1036768, 25'd4354425}, '{25'd2695596, -25'd414707, 25'd3939718, 25'd3317657, -25'd1368534, 25'd663531, -25'd2902950, -25'd1327063, -25'd1866182}, '{-25'd2239418, 25'd2737067, -25'd3193245, 25'd663531, -25'd207354, 25'd1824711, -25'd3981188, -25'd2861479, 25'd331766}, '{25'd4769132, 25'd2405301, -25'd2985891, 25'd1741770, 25'd1285592, -25'd2280889, -25'd3649423, 25'd539119, -25'd1078239}}},
    '{'{'{-25'd1800344, -25'd180034, 25'd2220425, -25'd2040390, -25'd2400459, -25'd1860356, 25'd0, 25'd3360643, -25'd1860356}, '{-25'd2820539, 25'd1020195, -25'd1980379, -25'd2880551, 25'd5281010, 25'd1020195, -25'd2520482, 25'd3720711, 25'd3480666}, '{25'd4200803, 25'd3600689, 25'd3300631, -25'd2160413, 25'd1800344, -25'd960184, 25'd2580493, 25'd1080207, -25'd1800344}, '{25'd4020769, 25'd3240620, 25'd2700516, 25'd360069, -25'd1860356, 25'd60011, 25'd960184, -25'd4080780, 25'd780149}, '{-25'd1620310, -25'd2700516, 25'd3960757, 25'd1860356, 25'd3780723, 25'd3060585, -25'd960184, 25'd5100975, 25'd5521056}, '{25'd3720711, 25'd4080780, 25'd6241193, 25'd4740907, 25'd7141366, 25'd7441423, 25'd4980952, 25'd2760528, -25'd1680321}, '{25'd2040390, -25'd1800344, -25'd120023, 25'd240046, 25'd7621457, 25'd7141366, 25'd3660700, 25'd2580493, 25'd4200803}, '{-25'd720138, 25'd4260815, 25'd4680895, -25'd2400459, 25'd1020195, 25'd2820539, 25'd2400459, 25'd2400459, 25'd4800918}, '{25'd4620884, -25'd2220425, -25'd1380264, -25'd2460470, -25'd960184, 25'd3840734, -25'd1800344, -25'd120023, -25'd1860356}}, '{'{25'd2880551, 25'd1620310, -25'd1560298, 25'd3960757, 25'd4860930, -25'd4320826, 25'd3960757, 25'd1920367, -25'd5401033}, '{25'd3360643, -25'd2820539, 25'd2940562, -25'd1500287, 25'd1140218, 25'd2580493, 25'd720138, -25'd780149, 25'd1440275}, '{-25'd1980379, 25'd2940562, -25'd2640505, -25'd4980952, -25'd480092, -25'd3420654, -25'd4500861, -25'd2760528, -25'd2280436}, '{-25'd5641079, -25'd360069, -25'd1080207, 25'd600115, 25'd2580493, -25'd1680321, -25'd3900746, -25'd2940562, -25'd3960757}, '{-25'd120023, 25'd600115, 25'd3060585, 25'd420080, -25'd2400459, -25'd2580493, 25'd5461044, 25'd3360643, -25'd1260241}, '{-25'd3540677, 25'd3960757, -25'd420080, 25'd2580493, -25'd1980379, -25'd2520482, 25'd3900746, 25'd2400459, 25'd3180608}, '{-25'd1500287, -25'd3900746, 25'd2520482, 25'd2400459, 25'd2340448, 25'd2940562, 25'd3120597, 25'd840161, -25'd4500861}, '{25'd240046, -25'd1740333, -25'd1740333, -25'd3720711, 25'd4500861, 25'd2760528, 25'd1560298, -25'd3300631, -25'd1860356}, '{25'd1860356, 25'd4020769, -25'd2160413, -25'd4740907, -25'd2100402, 25'd960184, -25'd5701090, -25'd2160413, -25'd5701090}}, '{'{25'd3240620, -25'd2940562, -25'd600115, -25'd540103, -25'd4200803, -25'd2760528, -25'd180034, 25'd1920367, 25'd720138}, '{-25'd2700516, 25'd4200803, -25'd1020195, -25'd2640505, -25'd4080780, 25'd1260241, -25'd1860356, -25'd1020195, -25'd3720711}, '{25'd3300631, -25'd2160413, -25'd3840734, -25'd4860930, -25'd5220998, -25'd2460470, -25'd1020195, 25'd3000574, 25'd900172}, '{-25'd2160413, -25'd4380838, 25'd60011, -25'd2220425, -25'd4440849, 25'd3720711, 25'd60011, -25'd4800918, -25'd900172}, '{-25'd300057, -25'd4620884, -25'd3600689, 25'd4380838, 25'd1500287, 25'd780149, -25'd4140792, 25'd0, -25'd240046}, '{25'd840161, 25'd4260815, -25'd900172, -25'd2520482, -25'd960184, -25'd420080, -25'd3000574, -25'd1080207, 25'd3000574}, '{-25'd5160987, 25'd2400459, -25'd4260815, 25'd1920367, -25'd1380264, 25'd120023, -25'd960184, -25'd720138, -25'd180034}, '{-25'd2220425, 25'd660126, -25'd3540677, 25'd3660700, 25'd2580493, 25'd4020769, 25'd2700516, -25'd2340448, -25'd3780723}, '{25'd1200230, 25'd720138, -25'd2760528, 25'd3000574, -25'd4620884, -25'd300057, 25'd2940562, -25'd5401033, 25'd1920367}}},
    '{'{'{-25'd2845757, 25'd3492521, -25'd86235, -25'd1810937, -25'd4397989, 25'd2112759, 25'd2543935, -25'd1854054, 25'd4699812}, '{-25'd3492521, 25'd344940, 25'd3276933, -25'd1983407, 25'd4570459, -25'd1164174, 25'd86235, -25'd43118, 25'd4311754}, '{25'd1810937, 25'd3492521, 25'd2845757, 25'd3578756, 25'd905468, -25'd862351, 25'd4484224, -25'd2888875, -25'd1681584}, '{-25'd172470, 25'd2371465, 25'd2069642, 25'd2845757, 25'd1810937, -25'd3104463, 25'd1250409, -25'd1638466, -25'd4441106}, '{-25'd4009931, 25'd1810937, -25'd1336644, 25'd4139284, 25'd732998, 25'd905468, -25'd4182401, 25'd129353, -25'd646763}, '{25'd1854054, -25'd1077938, 25'd3837461, 25'd732998, -25'd4786047, -25'd2802640, -25'd3751226, -25'd2414582, -25'd689881}, '{25'd2069642, -25'd2328347, 25'd4354871, -25'd2457700, 25'd43118, 25'd1379761, 25'd0, -25'd215588, 25'd4397989}, '{-25'd474293, 25'd4311754, 25'd4441106, -25'd2802640, -25'd4354871, -25'd1681584, 25'd3837461, -25'd2069642, -25'd3664991}, '{25'd474293, 25'd2026524, -25'd4053049, 25'd1121056, -25'd2802640, 25'd3664991, -25'd3837461, -25'd2026524, -25'd1595349}}, '{'{25'd1509114, 25'd4268636, 25'd3233815, -25'd1164174, -25'd1681584, 25'd3233815, -25'd3018228, 25'd5475927, -25'd1638466}, '{25'd732998, -25'd5130987, 25'd1983407, 25'd2673287, -25'd819233, -25'd3147580, -25'd2457700, -25'd732998, 25'd948586}, '{-25'd1638466, -25'd2112759, 25'd862351, -25'd689881, -25'd3147580, 25'd3147580, 25'd3708108, -25'd2026524, -25'd43118}, '{-25'd2845757, -25'd4397989, -25'd2587052, -25'd1121056, 25'd86235, -25'd4311754, 25'd2716405, 25'd86235, -25'd1034821}, '{25'd1681584, -25'd3061345, -25'd4699812, -25'd5519045, -25'd4742929, -25'd2975110, -25'd3621873, -25'd431175, 25'd4570459}, '{-25'd1810937, 25'd2242112, 25'd2371465, -25'd1077938, 25'd3104463, -25'd86235, -25'd2371465, -25'd2802640, -25'd3363168}, '{25'd2630170, -25'd3061345, -25'd3406285, 25'd86235, -25'd517410, -25'd4570459, -25'd3233815, 25'd4829164, -25'd3794343}, '{-25'd1681584, -25'd2285229, -25'd1897172, -25'd3535638, -25'd3363168, 25'd4182401, -25'd3578756, -25'd689881, -25'd129353}, '{25'd215588, 25'd431175, -25'd3233815, -25'd3578756, -25'd3664991, 25'd3578756, 25'd1293526, 25'd560528, 25'd1379761}}, '{'{25'd1207291, -25'd603646, 25'd3104463, 25'd5087869, 25'd1854054, 25'd1207291, -25'd1681584, -25'd819233, -25'd991703}, '{25'd646763, 25'd3449403, 25'd3104463, 25'd1121056, 25'd1034821, -25'd2543935, 25'd4053049, -25'd258705, -25'd4182401}, '{25'd3406285, -25'd2673287, -25'd2759522, -25'd4786047, 25'd1293526, 25'd4182401, 25'd3406285, 25'd2543935, -25'd3621873}, '{-25'd3966813, 25'd2543935, -25'd689881, 25'd3147580, 25'd1465996, 25'd3449403, -25'd3449403, -25'd1121056, 25'd301823}, '{-25'd1810937, 25'd4354871, -25'd2587052, 25'd3492521, -25'd2975110, -25'd2630170, -25'd5174105, 25'd3708108, -25'd1121056}, '{-25'd4009931, -25'd1638466, 25'd1422879, -25'd2888875, 25'd3708108, 25'd1681584, -25'd301823, 25'd431175, 25'd2285229}, '{25'd4009931, 25'd1767819, -25'd2543935, -25'd4009931, -25'd172470, 25'd3147580, -25'd603646, 25'd2543935, 25'd4053049}, '{-25'd4699812, 25'd388058, 25'd2630170, -25'd3966813, 25'd4268636, 25'd3018228, 25'd3233815, -25'd862351, -25'd1422879}, '{-25'd4915399, 25'd3147580, 25'd2457700, 25'd4786047, 25'd4182401, -25'd129353, -25'd2328347, 25'd2328347, 25'd4570459}}},
    '{'{'{25'd3678105, -25'd720453, -25'd1971767, 25'd3829779, -25'd4512314, 25'd606698, 25'd3109326, -25'd2047605, -25'd568779}, '{-25'd2085523, -25'd2275116, 25'd947965, 25'd3450593, 25'd1971767, -25'd1099640, 25'd3298919, 25'd1782174, 25'd2085523}, '{-25'd2275116, -25'd3261000, -25'd3640186, 25'd417105, -25'd4019372, 25'd4246884, -25'd4133128, -25'd758372, 25'd2692221}, '{-25'd1820093, 25'd379186, 25'd910046, -25'd2085523, -25'd2275116, -25'd2692221, -25'd4360639, 25'd4777744, -25'd1365070}, '{-25'd3753942, -25'd3905616, -25'd3223081, 25'd2730139, -25'd985884, -25'd3640186, -25'd644616, -25'd2426791, -25'd4133128}, '{-25'd2388872, -25'd2047605, 25'd189593, -25'd4588151, -25'd2123442, 25'd1744256, -25'd2464709, -25'd720453, -25'd1440907}, '{25'd1820093, -25'd1023802, -25'd1327151, 25'd4284802, -25'd1858012, -25'd4284802, -25'd3261000, 25'd4626070, -25'd2199279}, '{25'd2237198, -25'd2957651, 25'd417105, -25'd3261000, -25'd113756, -25'd113756, 25'd2388872, 25'd4398558, -25'd3602267}, '{-25'd568779, -25'd1933849, 25'd3374756, -25'd4512314, 25'd3867698, 25'd379186, -25'd2805977, -25'd1137558, 25'd3412674}}, '{'{-25'd4739825, -25'd682535, -25'd2199279, -25'd1137558, -25'd2464709, -25'd2730139, -25'd4626070, -25'd3450593, -25'd455023}, '{-25'd4057291, 25'd3678105, -25'd3298919, 25'd4701907, -25'd4095209, -25'd1895930, 25'd1554663, -25'd2995570, -25'd3602267}, '{25'd1213395, 25'd3185163, -25'd1933849, -25'd379186, -25'd2692221, -25'd3185163, -25'd530860, 25'd4701907, 25'd1706337}, '{-25'd1592581, 25'd2730139, 25'd1554663, 25'd1933849, -25'd151674, 25'd1478826, -25'd4019372, -25'd1175477, -25'd4739825}, '{-25'd1592581, 25'd4588151, 25'd2199279, -25'd265430, 25'd606698, -25'd2161360, -25'd1289233, -25'd3526430, -25'd303349}, '{25'd1630500, 25'd1402988, 25'd3109326, -25'd3261000, -25'd2692221, -25'd4322721, 25'd910046, -25'd1402988, -25'd4550232}, '{-25'd1440907, 25'd2426791, 25'd3753942, -25'd1630500, 25'd2881814, 25'd227512, -25'd2805977, -25'd3943535, 25'd682535}, '{25'd2919732, -25'd3261000, 25'd1516744, 25'd4436477, -25'd3867698, 25'd2957651, 25'd1706337, 25'd4095209, 25'd910046}, '{25'd2161360, 25'd2768058, -25'd1213395, -25'd4322721, 25'd0, -25'd2313035, -25'd2730139, -25'd265430, -25'd1061721}}, '{'{25'd2843895, -25'd3829779, 25'd4588151, -25'd3185163, 25'd1895930, 25'd1251314, 25'd1858012, -25'd1592581, 25'd1516744}, '{25'd4663988, 25'd4815663, -25'd4019372, -25'd3716023, -25'd4512314, -25'd3336837, 25'd2502628, -25'd1516744, -25'd4701907}, '{25'd1554663, -25'd1706337, 25'd2654302, 25'd872128, -25'd4057291, 25'd151674, 25'd4019372, -25'd3867698, -25'd4322721}, '{25'd1933849, -25'd37919, -25'd2350953, 25'd4246884, 25'd3791860, -25'd4588151, -25'd4512314, 25'd1782174, 25'd0}, '{25'd568779, -25'd1251314, 25'd1175477, 25'd4550232, -25'd1213395, -25'd303349, 25'd4663988, 25'd303349, -25'd189593}, '{25'd3071407, -25'd2654302, -25'd3981453, -25'd455023, 25'd4815663, 25'd3185163, -25'd3450593, 25'd37919, 25'd1023802}, '{-25'd227512, 25'd2919732, -25'd2730139, -25'd1365070, -25'd3298919, -25'd530860, -25'd3526430, 25'd492942, -25'd1820093}, '{-25'd1668419, 25'd2578465, -25'd2692221, 25'd0, -25'd3791860, -25'd1782174, -25'd3071407, -25'd910046, 25'd4436477}, '{25'd2237198, 25'd2275116, 25'd796291, -25'd1478826, -25'd985884, 25'd2843895, -25'd2199279, -25'd75837, 25'd1706337}}},
    '{'{'{-25'd4134743, 25'd2193945, -25'd1265738, -25'd1898607, 25'd4008170, -25'd4387891, -25'd2953388, -25'd1392312, -25'd4261317}, '{-25'd4092552, 25'd421913, -25'd3755022, 25'd1772033, 25'd928208, -25'd3544066, -25'd4387891, -25'd253148, 25'd4345700}, '{25'd3797213, -25'd3544066, -25'd2109563, 25'd4641038, -25'd1814224, 25'd3037771, -25'd1940798, 25'd4092552, 25'd4303508}, '{-25'd3628448, -25'd464104, -25'd3037771, 25'd3417492, 25'd3628448, 25'd1476694, -25'd3290918, 25'd1603268, -25'd464104}, '{25'd3164344, -25'd3797213, 25'd1772033, -25'd1307929, 25'd759443, 25'd5273907, 25'd5147334, -25'd1940798, 25'd3164344}, '{25'd2025180, -25'd3755022, -25'd3079962, 25'd970399, -25'd337530, -25'd632869, -25'd2320519, -25'd253148, -25'd1561077}, '{25'd4134743, 25'd2362710, 25'd4683230, -25'd4092552, 25'd1307929, -25'd3290918, 25'd1307929, 25'd4303508, 25'd2573667}, '{-25'd3839405, 25'd2911197, 25'd3248727, 25'd3375301, -25'd1603268, -25'd4387891, 25'd548486, -25'd2362710, -25'd843825}, '{25'd2911197, -25'd2869006, 25'd295339, -25'd2531475, 25'd1814224, -25'd2447093, 25'd2826814, -25'd2995579, -25'd548486}}, '{'{-25'd3459683, 25'd3839405, -25'd1181355, -25'd337530, 25'd337530, 25'd1012590, 25'd2995579, 25'd3417492, 25'd2109563}, '{25'd1223546, 25'd3670639, 25'd675060, 25'd84383, -25'd2700241, 25'd3206536, -25'd3839405, 25'd3333109, -25'd1687650}, '{-25'd3417492, -25'd1223546, -25'd3797213, -25'd2742432, 25'd2320519, -25'd379721, -25'd4387891, -25'd3965978, 25'd1814224}, '{25'd2742432, -25'd3755022, 25'd2911197, -25'd421913, 25'd337530, 25'd2362710, -25'd3797213, -25'd1096973, -25'd2784623}, '{-25'd1814224, 25'd4008170, 25'd3670639, 25'd295339, 25'd5020760, 25'd4978568, 25'd0, -25'd4134743, 25'd3375301}, '{25'd2700241, -25'd1012590, 25'd2362710, 25'd3459683, 25'd2700241, -25'd1603268, 25'd2911197, 25'd4387891, 25'd337530}, '{25'd2826814, -25'd1350120, 25'd4978568, -25'd4556656, 25'd1265738, -25'd3501874, -25'd2826814, 25'd1476694, -25'd2911197}, '{25'd3881596, -25'd632869, -25'd3544066, 25'd3459683, 25'd42191, 25'd4978568, 25'd3755022, -25'd2404902, -25'd3037771}, '{-25'd2193945, 25'd3712831, 25'd421913, -25'd4556656, -25'd3712831, -25'd1181355, 25'd675060, 25'd2995579, -25'd632869}}, '{'{25'd2826814, -25'd4345700, -25'd1434503, 25'd1096973, 25'd4387891, -25'd2869006, 25'd3459683, 25'd2278328, 25'd1561077}, '{25'd3164344, -25'd886016, -25'd2404902, 25'd632869, -25'd2869006, -25'd3839405, 25'd3670639, -25'd2236137, 25'd675060}, '{25'd3797213, 25'd2447093, -25'd2615858, -25'd1645459, -25'd2911197, -25'd717251, -25'd590678, 25'd2151754, -25'd421913}, '{-25'd4134743, -25'd717251, -25'd2067372, 25'd3586257, -25'd3164344, -25'd3670639, -25'd3923787, 25'd1392312, 25'd0}, '{-25'd886016, 25'd3037771, 25'd3501874, 25'd3712831, 25'd5358290, 25'd1561077, 25'd5062951, -25'd2911197, 25'd1518885}, '{25'd4345700, -25'd4261317, 25'd4809803, -25'd3670639, 25'd3037771, 25'd1012590, 25'd1350120, -25'd2151754, 25'd4851995}, '{-25'd4598847, 25'd4978568, 25'd2953388, -25'd3079962, 25'd886016, 25'd1096973, 25'd3417492, -25'd3670639, 25'd1603268}, '{25'd4936377, 25'd2742432, -25'd4092552, 25'd3755022, 25'd3501874, 25'd4725421, -25'd3839405, 25'd1181355, 25'd295339}, '{-25'd632869, 25'd4261317, -25'd2869006, 25'd506295, 25'd3544066, -25'd1476694, 25'd3333109, -25'd42191, 25'd1434503}}},
    '{'{'{25'd2303684, 25'd3602125, -25'd3853436, 25'd4649254, -25'd209426, 25'd1968603, -25'd4691139, -25'd2513110, -25'd2219914}, '{25'd4733024, -25'd2387455, 25'd2010488, 25'd837703, -25'd3979091, 25'd1633522, -25'd1089014, 25'd3392699, 25'd2848192}, '{-25'd3183273, 25'd1130900, 25'd83770, 25'd3350814, 25'd628278, -25'd3602125, -25'd2806306, -25'd125656, -25'd1172785}, '{25'd3099503, -25'd1549751, 25'd2596881, -25'd4942450, 25'd460737, -25'd1675407, 25'd3015732, 25'd1675407, 25'd3769665}, '{-25'd837703, -25'd1424096, -25'd3141388, -25'd3099503, -25'd251311, -25'd1424096, -25'd4774910, -25'd1842948, 25'd2638766}, '{25'd3979091, -25'd1424096, -25'd1172785, -25'd1759177, 25'd1005244, -25'd544507, 25'd3308929, -25'd2931962, -25'd4691139}, '{-25'd1465981, 25'd2387455, -25'd1675407, -25'd4900565, 25'd1382211, 25'd2010488, -25'd2513110, -25'd3727780, -25'd3811551}, '{-25'd2345570, 25'd3434584, -25'd837703, -25'd2052373, 25'd1633522, -25'd3602125, -25'd3015732, -25'd921474, -25'd1842948}, '{25'd4356058, 25'd586392, -25'd2178029, 25'd4607369, 25'd5235646, 25'd4356058, 25'd712048, 25'd4858680, 25'd1507866}}, '{'{-25'd4816795, 25'd544507, 25'd3350814, 25'd1214670, 25'd921474, 25'd4020976, 25'd2764421, 25'd2178029, 25'd2973847}, '{25'd3057618, 25'd4984335, 25'd2178029, -25'd2219914, 25'd3979091, -25'd3769665, 25'd963359, 25'd2554995, 25'd3141388}, '{-25'd3560240, 25'd1633522, 25'd1047129, 25'd4272288, -25'd167541, 25'd544507, -25'd1549751, -25'd2345570, -25'd3853436}, '{-25'd4439828, 25'd4104747, 25'd1842948, -25'd670163, -25'd1884833, -25'd4314173, -25'd837703, 25'd795818, 25'd3811551}, '{25'd586392, 25'd4607369, -25'd1340325, -25'd3811551, -25'd963359, -25'd418852, -25'd2596881, -25'd2931962, 25'd1675407}, '{-25'd2010488, -25'd5068106, -25'd4188517, 25'd1089014, -25'd3518354, 25'd2931962, -25'd712048, -25'd2052373, -25'd4649254}, '{25'd1089014, 25'd3602125, -25'd1884833, 25'd1382211, -25'd2345570, -25'd2806306, -25'd2052373, 25'd2471225, -25'd41885}, '{25'd2178029, 25'd3727780, -25'd2387455, -25'd3937206, -25'd4356058, 25'd3267043, -25'd1382211, -25'd2345570, -25'd4146632}, '{-25'd921474, 25'd167541, -25'd2596881, -25'd3979091, 25'd251311, 25'd3602125, -25'd2136144, 25'd2638766, -25'd1005244}}, '{'{25'd3350814, -25'd1005244, -25'd1801062, 25'd1130900, 25'd3350814, 25'd2973847, 25'd879589, -25'd1424096, 25'd1549751}, '{25'd41885, -25'd3685895, 25'd3602125, 25'd2806306, -25'd3937206, 25'd1759177, 25'd3769665, 25'd502622, 25'd2554995}, '{-25'd1256555, -25'd1214670, -25'd1465981, 25'd3350814, -25'd4774910, -25'd712048, 25'd2554995, -25'd4523599, 25'd2387455}, '{-25'd3937206, 25'd4607369, 25'd4272288, 25'd2010488, 25'd4146632, -25'd4104747, 25'd586392, -25'd4356058, 25'd1298440}, '{-25'd1842948, 25'd3979091, 25'd293196, -25'd3895321, 25'd3727780, 25'd1214670, -25'd4858680, 25'd1382211, 25'd879589}, '{-25'd2052373, 25'd2890077, -25'd209426, -25'd5319417, -25'd4774910, 25'd1759177, 25'd3267043, 25'd4020976, 25'd2554995}, '{25'd1298440, -25'd921474, -25'd3099503, -25'd1549751, -25'd3392699, 25'd4523599, -25'd83770, 25'd1884833, 25'd1424096}, '{25'd209426, -25'd2345570, 25'd2387455, 25'd1005244, -25'd2680651, 25'd4523599, -25'd921474, -25'd2219914, -25'd4020976}, '{25'd3015732, -25'd1549751, -25'd1591637, 25'd5319417, -25'd712048, 25'd251311, 25'd3015732, -25'd1340325, 25'd3560240}}},
    '{'{'{25'd1699936, 25'd2174337, 25'd1739469, 25'd2609204, -25'd1502269, -25'd118600, -25'd1699936, 25'd4823074, 25'd2174337}, '{-25'd4664941, 25'd3281272, 25'd711601, 25'd948802, -25'd948802, -25'd4783541, -25'd1027868, 25'd1067402, -25'd1383669}, '{-25'd4071940, 25'd2213870, 25'd830201, -25'd316267, 25'd276734, 25'd434867, 25'd4348674, -25'd4862608, 25'd79067}, '{25'd1146468, -25'd513934, -25'd790668, 25'd1779003, 25'd355801, 25'd4190540, 25'd118600, 25'd4704474, -25'd3281272}, '{-25'd3992873, 25'd3676606, 25'd4230073, 25'd1344135, -25'd3478939, 25'd2767338, -25'd4427740, -25'd1620869, 25'd4783541}, '{25'd1067402, 25'd434867, -25'd2727804, 25'd197667, -25'd1699936, 25'd3399872, -25'd1186002, -25'd1660403, 25'd4506807}, '{25'd2134803, -25'd3834739, -25'd3004538, -25'd3716139, 25'd3716139, -25'd4071940, -25'd39533, -25'd830201, 25'd355801}, '{25'd4111473, -25'd2095270, 25'd1660403, 25'd39533, 25'd2332470, 25'd4388207, 25'd276734, -25'd4190540, 25'd1660403}, '{-25'd790668, 25'd1383669, 25'd2332470, -25'd2411537, 25'd3320805, 25'd3637072, -25'd39533, 25'd3399872, 25'd1106935}}, '{'{25'd3992873, 25'd2846405, 25'd2569671, 25'd3992873, -25'd4585874, 25'd948802, 25'd4704474, -25'd2530137, 25'd355801}, '{25'd237200, -25'd2925471, -25'd1383669, -25'd434867, 25'd4032406, 25'd3637072, -25'd1146468, -25'd1344135, 25'd1265069}, '{25'd276734, -25'd1858070, 25'd2648738, 25'd3241738, 25'd830201, 25'd1502269, -25'd3241738, 25'd2648738, 25'd2174337}, '{-25'd1541802, -25'd553468, -25'd434867, -25'd3044071, -25'd3795206, -25'd4506807, 25'd2372004, -25'd909268, -25'd2016203}, '{-25'd1581336, -25'd158134, 25'd4902141, -25'd5060275, -25'd1344135, -25'd790668, 25'd1937136, 25'd2095270, -25'd3755673}, '{25'd1225535, 25'd3004538, 25'd1344135, 25'd2332470, 25'd3795206, 25'd2530137, -25'd2648738, -25'd1186002, -25'd3992873}, '{25'd4546341, 25'd5020741, 25'd1462736, -25'd2965005, 25'd1225535, 25'd4744008, 25'd3439405, 25'd4862608, -25'd1541802}, '{25'd1502269, -25'd1541802, 25'd3162672, -25'd513934, -25'd3716139, 25'd1858070, 25'd909268, 25'd1383669, 25'd3795206}, '{-25'd2609204, 25'd2965005, 25'd2569671, -25'd2965005, -25'd4506807, -25'd3044071, 25'd3676606, 25'd553468, -25'd1106935}}, '{'{-25'd3439405, 25'd2846405, -25'd3399872, -25'd553468, 25'd3874273, 25'd4467274, 25'd79067, -25'd2372004, -25'd3439405}, '{-25'd1897603, 25'd2688271, 25'd4071940, -25'd4388207, -25'd3874273, -25'd988335, 25'd2490604, 25'd3795206, 25'd4388207}, '{-25'd2411537, -25'd276734, 25'd4388207, 25'd3162672, 25'd1067402, 25'd2411537, -25'd2806871, -25'd988335, -25'd1423202}, '{-25'd3004538, 25'd1067402, 25'd237200, -25'd869735, 25'd2095270, -25'd2688271, 25'd751135, 25'd4585874, -25'd2569671}, '{25'd4546341, -25'd3004538, -25'd948802, 25'd513934, -25'd2609204, 25'd2925471, -25'd4744008, 25'd4071940, -25'd1344135}, '{25'd355801, -25'd1383669, 25'd3676606, -25'd4783541, -25'd1620869, -25'd1739469, -25'd1858070, -25'd1383669, 25'd2332470}, '{25'd3083605, -25'd1858070, -25'd4704474, 25'd3360339, -25'd3478939, -25'd2925471, 25'd1186002, -25'd2411537, 25'd4071940}, '{-25'd3123138, 25'd4506807, 25'd1067402, 25'd1779003, -25'd1937136, -25'd1067402, -25'd3913806, -25'd1186002, 25'd1581336}, '{-25'd434867, -25'd2292937, 25'd2411537, 25'd3953340, -25'd4190540, -25'd3123138, -25'd3518472, -25'd3162672, -25'd3360339}}},
    '{'{'{25'd164581, 25'd4649427, 25'd41145, -25'd2921321, -25'd740617, 25'd3456211, -25'd3785374, 25'd2345286, 25'd946344}, '{-25'd2921321, -25'd3373920, 25'd3703083, 25'd2427577, 25'd452599, 25'd1974978, 25'd2221850, -25'd1522379, -25'd740617}, '{-25'd3703083, 25'd2221850, -25'd164581, -25'd4402555, -25'd4525991, -25'd617181, 25'd1686960, 25'd2921321, 25'd452599}, '{25'd3579647, 25'd246872, -25'd699471, 25'd2180705, 25'd2139559, 25'd4608281, 25'd4155682, 25'd41145, -25'd4361409}, '{25'd4525991, 25'd2551013, 25'd2797885, 25'd4484845, 25'd1892687, 25'd2139559, 25'd1522379, 25'd1481233, -25'd41145}, '{-25'd4279119, 25'd2509868, 25'd205727, -25'd3744229, 25'd1563524, 25'd3456211, 25'd1193216, 25'd4073392, 25'd2756740}, '{25'd3867665, 25'd781762, -25'd2633304, 25'd534890, -25'd3579647, -25'd2468722, 25'd1522379, -25'd4937444, 25'd3415066}, '{25'd2509868, -25'd4649427, -25'd740617, 25'd329163, 25'd3661938, 25'd1892687, 25'd1152070, -25'd1563524, 25'd2509868}, '{-25'd2057269, -25'd1234361, -25'd905198, 25'd3044757, -25'd699471, 25'd3209339, -25'd1522379, -25'd1522379, -25'd3373920}}, '{'{-25'd1316652, -25'd4237973, 25'd2509868, -25'd1974978, -25'd2468722, -25'd1810396, 25'd1481233, 25'd4155682, 25'd2839031}, '{25'd4608281, 25'd2921321, 25'd4155682, -25'd2221850, 25'd3949956, -25'd3127048, 25'd3497356, -25'd822907, 25'd658326}, '{-25'd2345286, 25'd1769251, 25'd864053, -25'd2262995, 25'd2962467, -25'd4814008, -25'd3291630, 25'd411454, 25'd4402555}, '{-25'd123436, 25'd2797885, -25'd2386431, 25'd2386431, -25'd4402555, 25'd2880176, 25'd1316652, 25'd4567136, 25'd2016123}, '{25'd2221850, 25'd781762, 25'd1645815, -25'd2057269, -25'd905198, -25'd5266607, -25'd5019735, 25'd2098414, 25'd3620793}, '{25'd4279119, -25'd946344, -25'd2345286, 25'd82291, 25'd2633304, -25'd2715594, -25'd493744, 25'd2427577, -25'd4937444}, '{25'd1275506, -25'd411454, 25'd2756740, 25'd2880176, -25'd3044757, -25'd4731718, -25'd905198, -25'd1275506, -25'd2674449}, '{-25'd164581, -25'd4690572, 25'd4484845, -25'd1810396, 25'd1028634, -25'd2057269, -25'd3127048, 25'd82291, -25'd3949956}, '{25'd2839031, -25'd164581, -25'd1810396, -25'd4279119, -25'd3579647, 25'd3497356, 25'd2098414, -25'd4361409, -25'd4690572}}, '{'{-25'd4649427, -25'd205727, -25'd5266607, 25'd3291630, -25'd4608281, 25'd822907, 25'd2427577, -25'd4155682, -25'd5102026}, '{-25'd4361409, -25'd1810396, -25'd3003612, -25'd1481233, 25'd1316652, -25'd2139559, 25'd493744, -25'd5019735, -25'd4402555}, '{-25'd4196828, 25'd2016123, 25'd1563524, 25'd2633304, -25'd452599, 25'd1769251, -25'd1275506, -25'd3332775, -25'd3085903}, '{-25'd205727, 25'd576035, 25'd2797885, -25'd370308, 25'd1440088, 25'd4196828, 25'd2921321, -25'd1933832, 25'd3044757}, '{-25'd493744, -25'd4608281, 25'd3209339, -25'd4772863, -25'd3908810, 25'd3579647, -25'd4690572, -25'd2715594, -25'd4361409}, '{-25'd3291630, -25'd740617, -25'd946344, -25'd4484845, 25'd1357797, 25'd2797885, -25'd2139559, 25'd370308, 25'd2345286}, '{-25'd4567136, -25'd3415066, 25'd2715594, 25'd3332775, -25'd2180705, -25'd3497356, -25'd905198, -25'd2962467, 25'd205727}, '{-25'd4114537, 25'd3456211, -25'd4525991, 25'd3497356, 25'd2797885, 25'd987489, 25'd2180705, 25'd2674449, -25'd3497356}, '{25'd3415066, 25'd1152070, 25'd2098414, 25'd452599, -25'd3456211, -25'd4855154, -25'd2427577, 25'd822907, 25'd534890}}},
    '{'{'{-25'd582290, 25'd3909662, -25'd3119411, -25'd4866282, -25'd1830055, -25'd5199019, 25'd2121200, 25'd3119411, -25'd3992846}, '{-25'd956619, -25'd2121200, -25'd1663686, -25'd3161003, -25'd1497317, 25'd1663686, -25'd1497317, -25'd5323795, 25'd4200807}, '{25'd1414133, -25'd2204384, -25'd83184, -25'd3784886, -25'd4991058, 25'd2953043, 25'd2661898, -25'd2703490, 25'd3119411}, '{25'd1538910, 25'd4450360, -25'd4408768, 25'd3368964, 25'd998212, -25'd1206172, -25'd1913239, 25'd3826478, -25'd1830055}, '{25'd790251, -25'd915027, 25'd665474, 25'd2911450, -25'd1746870, -25'd3951254, -25'd4450360, -25'd3202596, 25'd1788462}, '{25'd2869858, 25'd83184, -25'd457514, 25'd1039804, 25'd2287568, 25'd374329, -25'd3951254, 25'd249553, 25'd1622094}, '{25'd3743293, -25'd4783097, -25'd1122988, 25'd2869858, -25'd915027, -25'd5199019, -25'd1622094, -25'd1788462, 25'd3244188}, '{25'd2745082, -25'd5032650, 25'd831843, -25'd3493741, 25'd1164580, 25'd3452148, -25'd873435, -25'd1663686, 25'd915027}, '{-25'd3410556, -25'd3410556, -25'd873435, 25'd2245976, -25'd1455725, 25'd1372541, 25'd4949466, -25'd3535333, -25'd4450360}}, '{'{25'd956619, 25'd2079607, -25'd582290, 25'd1705278, 25'd540698, 25'd249553, 25'd2162792, 25'd4076031, -25'd2869858}, '{25'd2370753, 25'd956619, 25'd3285780, -25'd5074242, 25'd3161003, 25'd3743293, -25'd2038015, 25'd1039804, 25'd2911450}, '{25'd3368964, -25'd3826478, 25'd166369, -25'd291145, -25'd1372541, -25'd3701701, 25'd1788462, 25'd3784886, 25'd790251}, '{-25'd956619, -25'd540698, 25'd3119411, -25'd3784886, 25'd3660109, 25'd207961, 25'd623882, -25'd3452148, -25'd5115834}, '{25'd1538910, -25'd1164580, -25'd3660109, 25'd3618517, -25'd41592, 25'd2953043, -25'd207961, -25'd1039804, -25'd41592}, '{-25'd2204384, -25'd457514, 25'd1746870, -25'd207961, 25'd2537121, 25'd2329160, -25'd166369, -25'd1663686, 25'd415921}, '{25'd457514, -25'd582290, -25'd2953043, 25'd4450360, 25'd4117623, -25'd332737, 25'd3743293, 25'd1705278, 25'd1497317}, '{25'd3327372, 25'd3826478, 25'd1206172, 25'd4533544, -25'd1871647, 25'd1039804, 25'd1081396, -25'd3701701, -25'd3452148}, '{-25'd998212, 25'd3161003, -25'd2121200, -25'd2162792, 25'd2204384, -25'd1247764, 25'd956619, 25'd1372541, -25'd1705278}}, '{'{-25'd5074242, 25'd3618517, 25'd457514, -25'd4283991, 25'd1497317, 25'd3743293, -25'd3036227, 25'd2495529, -25'd3951254}, '{25'd2911450, -25'd1206172, 25'd1081396, -25'd2828266, 25'd2370753, -25'd166369, -25'd3909662, -25'd4783097, 25'd4325584}, '{-25'd4616729, 25'd1372541, 25'd3285780, 25'd540698, 25'd707067, 25'd4533544, 25'd1414133, -25'd3410556, 25'd457514}, '{25'd1663686, -25'd4242399, 25'd4783097, 25'd3452148, 25'd2745082, -25'd3077819, 25'd3368964, 25'd3493741, 25'd207961}, '{-25'd3493741, -25'd4283991, 25'd1330949, -25'd374329, -25'd1039804, 25'd3368964, 25'd2537121, -25'd1580502, -25'd2828266}, '{-25'd1996423, -25'd3868070, 25'd2412345, 25'd0, 25'd790251, -25'd2578713, 25'd415921, -25'd3660109, -25'd4283991}, '{-25'd2370753, -25'd4824689, -25'd707067, -25'd3368964, -25'd332737, -25'd2079607, 25'd2412345, -25'd1746870, -25'd2537121}, '{-25'd1122988, 25'd1247764, 25'd4907874, 25'd4866282, 25'd1247764, -25'd3161003, 25'd4159215, -25'd582290, -25'd3202596}, '{25'd4242399, 25'd2620305, 25'd1330949, 25'd4907874, -25'd2786674, 25'd3618517, -25'd2079607, -25'd4367176, 25'd3576925}}},
    '{'{'{25'd702947, 25'd3676955, 25'd3785101, 25'd1514040, 25'd4001392, 25'd1189603, 25'd162219, 25'd4812485, -25'd4433975}, '{25'd2433279, -25'd2865862, 25'd5028777, -25'd54073, 25'd5299141, 25'd2974008, 25'd3136226, -25'd3460664, 25'd162219}, '{25'd4109538, -25'd2000696, -25'd324437, -25'd3406591, -25'd1838478, -25'd919239, -25'd1676259, 25'd5136923, -25'd4163611}, '{25'd1838478, -25'd1622186, -25'd3406591, -25'd1730332, 25'd2000696, 25'd1892550, 25'd0, -25'd3460664, 25'd4650267}, '{-25'd3136226, 25'd3028081, 25'd5136923, 25'd757020, 25'd5082850, 25'd3244372, 25'd973312, -25'd2974008, 25'd5082850}, '{-25'd2919935, -25'd324437, 25'd4920631, -25'd1946623, 25'd3244372, 25'd486656, 25'd3514736, 25'd4542121, 25'd1676259}, '{-25'd4001392, -25'd6650963, 25'd919239, -25'd3785101, 25'd2541425, 25'd2595498, -25'd594802, -25'd4001392, -25'd486656}, '{-25'd3514736, 25'd2379206, 25'd1730332, -25'd3136226, -25'd1243676, -25'd4217684, -25'd4596194, -25'd216291, -25'd1784405}, '{25'd1838478, -25'd1946623, 25'd324437, 25'd1838478, -25'd3622882, 25'd540729, -25'd5461360, -25'd4433975, -25'd3893247}}, '{'{-25'd54073, -25'd3839174, -25'd2649571, 25'd3731028, -25'd5082850, 25'd702947, 25'd1135530, -25'd4379902, 25'd378510}, '{25'd4217684, -25'd3352518, 25'd2919935, -25'd1730332, -25'd811093, -25'd1676259, 25'd2919935, 25'd2108842, -25'd1730332}, '{-25'd1568113, -25'd919239, 25'd4217684, 25'd3731028, 25'd3731028, -25'd540729, 25'd432583, 25'd1892550, -25'd1622186}, '{-25'd3244372, -25'd540729, 25'd3568809, 25'd3082154, -25'd1676259, -25'd1297749, -25'd4055465, -25'd108146, -25'd2433279}, '{25'd54073, -25'd757020, -25'd2865862, -25'd3514736, -25'd540729, -25'd1676259, 25'd1243676, -25'd2325133, -25'd2919935}, '{-25'd2487352, 25'd3082154, -25'd1946623, 25'd3406591, 25'd648874, 25'd4704340, 25'd2325133, 25'd4812485, 25'd811093}, '{-25'd2216988, 25'd3028081, -25'd757020, 25'd3136226, 25'd2703643, -25'd3406591, -25'd2433279, 25'd648874, -25'd6434671}, '{-25'd6921327, -25'd6272453, 25'd702947, -25'd2000696, -25'd324437, -25'd1243676, 25'd2487352, -25'd1459967, -25'd4271757}, '{-25'd2379206, 25'd2216988, 25'd2649571, 25'd1730332, 25'd1730332, -25'd3568809, -25'd702947, -25'd4974704, 25'd757020}}, '{'{-25'd757020, 25'd4055465, -25'd5190995, -25'd2108842, -25'd1189603, -25'd3514736, -25'd1135530, 25'd486656, 25'd2379206}, '{-25'd4217684, -25'd4217684, -25'd3514736, -25'd1892550, -25'd3947319, -25'd2919935, 25'd2216988, 25'd2865862, 25'd2865862}, '{25'd324437, -25'd4271757, 25'd1838478, 25'd2000696, 25'd1784405, -25'd4433975, -25'd5407287, -25'd5948016, -25'd2271060}, '{25'd54073, -25'd811093, -25'd4433975, 25'd2000696, -25'd1676259, 25'd0, 25'd2649571, 25'd973312, -25'd3460664}, '{-25'd2649571, 25'd108146, -25'd54073, 25'd2811789, 25'd3298445, -25'd2974008, -25'd1351822, 25'd2757716, -25'd3352518}, '{25'd1784405, -25'd3622882, 25'd2433279, 25'd2541425, 25'd2919935, -25'd270364, -25'd1297749, 25'd3785101, -25'd1622186}, '{-25'd5569506, 25'd973312, -25'd2487352, 25'd3460664, -25'd2162915, -25'd1135530, -25'd3028081, -25'd3244372, -25'd1027385}, '{-25'd6110234, -25'd1946623, 25'd973312, -25'd4920631, 25'd1730332, -25'd270364, -25'd5839870, -25'd4866558, -25'd1784405}, '{-25'd5245068, 25'd216291, -25'd919239, -25'd540729, 25'd54073, 25'd1189603, -25'd5785797, -25'd162219, 25'd3676955}}},
    '{'{'{-25'd1646596, 25'd3799837, 25'd2533224, 25'd1984359, -25'd126661, 25'd337763, -25'd3546514, 25'd4728685, -25'd2111020}, '{-25'd3166530, -25'd1266612, -25'd3588735, -25'd506645, 25'd1899918, -25'd2828767, 25'd3926498, 25'd84441, -25'd84441}, '{25'd1139951, 25'd4010939, -25'd1393273, -25'd3842057, 25'd2744326, 25'd3293192, -25'd2026579, 25'd886629, 25'd4095379}, '{25'd5361992, 25'd3039869, -25'd5277551, 25'd759967, -25'd1773257, -25'd4475363, 25'd2068800, 25'd2617665, -25'd2828767}, '{-25'd211102, -25'd1688816, -25'd5193110, -25'd464424, 25'd2364343, -25'd3166530, -25'd1731037, -25'd3462073, -25'd4475363}, '{25'd4897567, -25'd3293192, -25'd1477714, 25'd1182171, -25'd928849, 25'd2364343, -25'd928849, 25'd2702106, 25'd1224392}, '{25'd4897567, 25'd4728685, -25'd4095379, -25'd3757616, -25'd168882, -25'd379984, 25'd2702106, 25'd4095379, -25'd295543}, '{-25'd928849, 25'd3124310, 25'd802188, -25'd5319771, 25'd3208751, -25'd4686465, -25'd1182171, -25'd2997649, -25'd84441}, '{-25'd3630955, 25'd1731037, -25'd4939788, 25'd3208751, 25'd759967, 25'd3335412, -25'd295543, 25'd1773257, -25'd211102}}, '{'{-25'd3842057, -25'd84441, -25'd211102, 25'd464424, 25'd2786547, -25'd1308833, -25'd1688816, -25'd3588735, -25'd3757616}, '{25'd3166530, 25'd928849, 25'd2955428, -25'd4348702, 25'd2068800, 25'd253322, 25'd4053159, 25'd3208751, -25'd1899918}, '{-25'd1773257, -25'd1815477, 25'd3250971, 25'd1857698, 25'd3082090, -25'd971069, 25'd3546514, 25'd3462073, 25'd1308833}, '{25'd42220, -25'd3377632, -25'd1224392, -25'd3546514, -25'd4179820, 25'd1688816, 25'd3293192, 25'd2279902, -25'd2364343}, '{25'd4728685, 25'd4855347, -25'd4728685, -25'd5404212, -25'd3715396, -25'd2533224, -25'd2786547, 25'd802188, -25'd1984359}, '{25'd2448784, 25'd4813126, 25'd1984359, 25'd3419853, 25'd3377632, 25'd2406563, -25'd5319771, -25'd2491004, 25'd548865}, '{-25'd2406563, 25'd3968718, -25'd4390922, 25'd2153241, -25'd3293192, -25'd3293192, -25'd886629, -25'd844408, 25'd3250971}, '{25'd802188, -25'd1942139, 25'd3377632, 25'd3377632, -25'd2237682, 25'd4559804, -25'd886629, -25'd4306481, -25'd4137600}, '{25'd4010939, -25'd1393273, -25'd2913208, -25'd3377632, -25'd1393273, -25'd1731037, -25'd3504294, -25'd3082090, 25'd1055510}}, '{'{25'd675526, 25'd3926498, -25'd3842057, 25'd4095379, -25'd5277551, -25'd4010939, 25'd2111020, -25'd928849, 25'd3842057}, '{-25'd2870988, -25'd3419853, 25'd0, -25'd3082090, 25'd1013290, 25'd4348702, 25'd1688816, -25'd2068800, 25'd2617665}, '{-25'd1688816, -25'd1308833, 25'd1604375, -25'd3124310, -25'd4348702, -25'd1688816, -25'd2068800, 25'd3799837, 25'd3166530}, '{25'd717747, 25'd506645, 25'd844408, 25'd2153241, -25'd4264261, 25'd1519935, 25'd337763, 25'd295543, -25'd3799837}, '{25'd422204, -25'd3124310, -25'd2997649, -25'd4475363, 25'd253322, -25'd1435494, -25'd4179820, 25'd422204, 25'd42220}, '{25'd675526, -25'd548865, 25'd2913208, -25'd802188, 25'd3124310, 25'd1013290, -25'd591086, 25'd1266612, 25'd759967}, '{25'd4264261, 25'd0, 25'd422204, 25'd1519935, -25'd971069, -25'd3926498, 25'd2237682, 25'd3208751, 25'd2744326}, '{25'd2026579, 25'd4559804, 25'd1731037, 25'd2153241, -25'd379984, 25'd1731037, -25'd4264261, 25'd3462073, -25'd1773257}, '{25'd3419853, 25'd2111020, 25'd3968718, -25'd3335412, 25'd2237682, 25'd633306, 25'd1266612, 25'd1688816, 25'd3715396}}},
    '{'{'{-25'd2487149, -25'd5321342, -25'd2313627, 25'd57841, 25'd4164528, 25'd2602830, 25'd3123396, 25'd2313627, -25'd173522}, '{25'd1330335, 25'd1446017, -25'd4280210, -25'd4222369, 25'd5321342, 25'd4800776, -25'd3643962, 25'd1098973, -25'd2892034}, '{25'd2487149, -25'd1966583, -25'd2718512, -25'd2660671, 25'd636247, 25'd4106688, -25'd3354759, 25'd751929, -25'd4858616}, '{25'd520566, 25'd115681, 25'd1966583, -25'd1041132, 25'd3354759, 25'd6304633, 25'd4511572, -25'd3643962, -25'd751929}, '{25'd4858616, -25'd2487149, 25'd6362474, 25'd4453732, 25'd7287924, 25'd7345765, 25'd4916457, -25'd462725, -25'd3181237}, '{-25'd1908742, -25'd2255786, 25'd1272495, -25'd1793061, 25'd2602830, 25'd4164528, 25'd1850901, 25'd1503857, 25'd578407}, '{-25'd3239078, 25'd2082264, -25'd578407, 25'd3817484, 25'd2834193, 25'd4280210, 25'd2024423, -25'd404885, -25'd4106688}, '{-25'd3643962, 25'd2949874, -25'd4395891, 25'd2371467, 25'd1677379, 25'd2197945, 25'd289203, 25'd4800776, 25'd4106688}, '{-25'd5089979, 25'd1677379, -25'd1098973, -25'd578407, 25'd3239078, 25'd2949874, -25'd2487149, 25'd3875325, -25'd809769}}, '{'{25'd2834193, 25'd404885, 25'd983291, 25'd2602830, -25'd2255786, 25'd3239078, 25'd289203, -25'd3528281, -25'd2024423}, '{-25'd983291, 25'd1272495, 25'd3991006, -25'd3354759, 25'd3528281, 25'd5089979, -25'd231363, -25'd4916457, -25'd2024423}, '{-25'd520566, -25'd4395891, -25'd231363, -25'd2892034, -25'd1446017, 25'd4338050, 25'd3759644, -25'd4106688, -25'd1446017}, '{-25'd694088, 25'd578407, -25'd4280210, 25'd3123396, -25'd925451, -25'd2487149, 25'd3239078, -25'd2487149, -25'd5494864}, '{-25'd2602830, 25'd4974298, -25'd2487149, 25'd4627254, 25'd1388176, 25'd2660671, 25'd6767358, 25'd3759644, 25'd2082264}, '{25'd2197945, -25'd1272495, -25'd3528281, -25'd1793061, 25'd5494864, 25'd4164528, -25'd1850901, -25'd2544990, 25'd4453732}, '{25'd1561698, 25'd3933166, 25'd3007715, 25'd5147820, 25'd1214654, 25'd2197945, 25'd1966583, 25'd4974298, -25'd751929}, '{25'd2892034, 25'd3239078, -25'd983291, -25'd578407, -25'd694088, 25'd1214654, 25'd2082264, -25'd4916457, -25'd3643962}, '{25'd2660671, -25'd5841908, 25'd2429308, -25'd4106688, 25'd694088, 25'd1272495, 25'd3701803, -25'd4048847, 25'd2255786}}, '{'{-25'd1156813, -25'd3412600, 25'd636247, -25'd6478155, -25'd3991006, 25'd1793061, 25'd1619539, -25'd1503857, 25'd2313627}, '{25'd1446017, -25'd1330335, -25'd1619539, -25'd5899748, 25'd1619539, -25'd173522, 25'd1388176, -25'd1388176, -25'd2429308}, '{-25'd404885, -25'd1677379, -25'd694088, -25'd3528281, 25'd4280210, -25'd925451, -25'd231363, 25'd3528281, 25'd3296918}, '{25'd520566, -25'd4222369, -25'd5552704, -25'd2776352, 25'd404885, -25'd809769, -25'd2429308, 25'd115681, -25'd5089979}, '{25'd1098973, -25'd231363, 25'd2313627, 25'd1214654, -25'd1156813, 25'd6651677, 25'd2082264, -25'd3759644, -25'd694088}, '{-25'd173522, -25'd3239078, 25'd2197945, -25'd3065556, 25'd173522, 25'd1272495, -25'd1561698, -25'd3991006, -25'd5205660}, '{-25'd2197945, -25'd2371467, 25'd925451, -25'd867610, 25'd4569413, -25'd3239078, -25'd3239078, -25'd2024423, 25'd3701803}, '{-25'd4974298, -25'd4280210, -25'd2776352, -25'd3759644, 25'd925451, 25'd3412600, 25'd462725, -25'd4106688, 25'd3817484}, '{25'd1619539, 25'd3123396, 25'd925451, -25'd4800776, -25'd1330335, 25'd809769, -25'd1908742, -25'd4453732, -25'd3123396}}},
    '{'{'{-25'd2576898, -25'd356801, -25'd237867, 25'd634313, -25'd4876283, 25'd4400548, -25'd4479837, -25'd3845524, -25'd2259741}, '{-25'd4241970, -25'd2378675, -25'd4717705, 25'd3250855, -25'd1625428, 25'd0, 25'd3766235, -25'd3845524, 25'd2061518}, '{25'd4400548, -25'd3250855, -25'd4162681, 25'd3369789, -25'd1823651, -25'd4321259, -25'd1387560, -25'd911825, 25'd832536}, '{25'd4876283, -25'd3686946, -25'd4202325, 25'd396446, 25'd1982229, -25'd3449078, 25'd673958, -25'd2537253, -25'd2418319}, '{-25'd2339030, -25'd2457964, 25'd3845524, 25'd158578, -25'd4717705, 25'd4400548, -25'd5034861, 25'd3686946, 25'd1149693}, '{25'd1070404, -25'd1506494, -25'd2497608, -25'd1982229, -25'd277512, -25'd3686946, 25'd4360903, 25'd2299385, 25'd4241970}, '{-25'd673958, -25'd3964458, -25'd4955572, 25'd3568012, -25'd158578, -25'd3568012, 25'd2220096, -25'd2259741, 25'd673958}, '{-25'd1823651, -25'd4836638, -25'd713602, 25'd3607657, -25'd3885169, 25'd1665072, 25'd713602, -25'd911825, -25'd79289}, '{-25'd2814765, -25'd277512, 25'd1982229, 25'd3131922, -25'd2576898, -25'd3211211, 25'd1466849, 25'd4360903, -25'd1863295}}, '{'{25'd4559126, -25'd158578, 25'd3211211, 25'd3369789, 25'd2656187, 25'd2854410, -25'd3369789, -25'd991114, -25'd475735}, '{25'd1347916, 25'd3488723, 25'd3369789, 25'd4241970, -25'd158578, 25'd1506494, 25'd1665072, -25'd3409434, -25'd4995217}, '{-25'd2061518, -25'd1387560, 25'd2378675, -25'd436090, -25'd4043747, 25'd3330144, 25'd2814765, 25'd317157, -25'd3092277}, '{-25'd872181, 25'd1070404, 25'd2894054, 25'd2220096, -25'd1744361, -25'd1030759, 25'd3409434, -25'd3449078, 25'd3409434}, '{-25'd1268626, -25'd1387560, -25'd4757349, -25'd713602, 25'd39645, -25'd1268626, -25'd4083391, -25'd2814765, -25'd2656187}, '{-25'd3369789, 25'd1823651, -25'd3290500, 25'd2061518, 25'd1506494, 25'd2101163, -25'd2457964, 25'd2973343, 25'd237867}, '{-25'd1744361, -25'd1546139, -25'd4083391, 25'd3726590, 25'd2775120, 25'd3250855, 25'd991114, -25'd4796994, 25'd3171566}, '{-25'd1189337, -25'd951470, 25'd1902940, 25'd1506494, -25'd4757349, 25'd2894054, -25'd2457964, -25'd1942584, 25'd555024}, '{25'd3805879, 25'd4241970, 25'd2735476, -25'd2695831, -25'd3607657, -25'd1704717, -25'd3924813, -25'd3211211, 25'd1308271}}, '{'{25'd3250855, -25'd3330144, -25'd3131922, -25'd713602, -25'd3528367, -25'd2497608, -25'd4559126, -25'd1982229, -25'd79289}, '{25'd1942584, -25'd3488723, 25'd1784006, 25'd4717705, 25'd4202325, 25'd2775120, -25'd2576898, 25'd1902940, -25'd198223}, '{-25'd753247, 25'd0, -25'd4638416, -25'd4519482, -25'd3845524, 25'd1665072, -25'd3726590, -25'd1308271, 25'd39645}, '{25'd3964458, -25'd2497608, -25'd1070404, -25'd1466849, -25'd3012988, -25'd2775120, -25'd2656187, -25'd1863295, -25'd673958}, '{25'd237867, 25'd4123036, 25'd3092277, -25'd872181, -25'd1070404, -25'd1744361, -25'd1704717, -25'd1585783, -25'd3766235}, '{-25'd1466849, -25'd3885169, -25'd634313, 25'd911825, 25'd79289, 25'd1665072, 25'd3250855, 25'd3845524, -25'd2259741}, '{25'd2021873, -25'd3250855, 25'd237867, 25'd2378675, 25'd3528367, -25'd3885169, -25'd1228982, 25'd3607657, -25'd4202325}, '{25'd2616542, 25'd1189337, -25'd4400548, 25'd872181, -25'd2299385, 25'd436090, -25'd4123036, 25'd1347916, -25'd4678060}, '{-25'd2656187, -25'd1070404, 25'd4440193, -25'd3250855, 25'd2537253, -25'd3211211, 25'd4400548, 25'd4440193, 25'd1942584}}},
    '{'{'{-25'd991646, -25'd3346806, 25'd4586364, -25'd1900655, -25'd2892301, 25'd2768346, 25'd4421089, -25'd826372, 25'd578460}, '{-25'd3759992, 25'd991646, -25'd3594718, 25'd991646, 25'd3553399, 25'd2355160, 25'd1611425, -25'd1652744, 25'd1446151}, '{-25'd1239558, 25'd1363514, -25'd2437797, 25'd2065930, -25'd1735381, -25'd3429443, 25'd2272523, 25'd4462408, 25'd5164824}, '{25'd661097, 25'd4792957, 25'd2107248, -25'd2974939, 25'd2189885, -25'd826372, -25'd1859337, 25'd5247461, 25'd4297134}, '{-25'd1652744, -25'd3553399, 25'd867690, 25'd123956, -25'd4503727, 25'd4545045, 25'd3264169, -25'd4007903, 25'd578460}, '{25'd1115602, 25'd4338452, -25'd1528788, -25'd1941974, -25'd2603071, -25'd3098894, 25'd4173178, 25'd2355160, -25'd3098894}, '{25'd3512080, 25'd2644390, 25'd330549, 25'd3016257, -25'd2561753, -25'd371867, -25'd3429443, 25'd41319, 25'd1735381}, '{-25'd867690, -25'd1074283, 25'd4669001, 25'd4421089, -25'd4462408, -25'd2355160, -25'd1694062, 25'd4834275, -25'd2727027}, '{25'd4007903, -25'd1652744, -25'd1652744, 25'd661097, -25'd537142, -25'd4131859, 25'd1570107, 25'd3305487, 25'd1239558}}, '{'{-25'd1694062, 25'd619779, -25'd3801311, -25'd4462408, -25'd2107248, -25'd991646, -25'd4462408, 25'd3512080, 25'd4503727}, '{25'd2396478, 25'd3305487, -25'd2603071, -25'd2272523, -25'd1735381, 25'd1156921, -25'd3140213, -25'd3057576, -25'd3677355}, '{-25'd3925266, -25'd661097, 25'd867690, 25'd3636036, 25'd2148567, -25'd4255815, -25'd4049222, -25'd4462408, 25'd1652744}, '{25'd3305487, 25'd3429443, 25'd3098894, 25'd5040868, 25'd1941974, 25'd619779, 25'd3181532, 25'd3512080, 25'd2561753}, '{25'd1611425, 25'd867690, -25'd4297134, 25'd2768346, -25'd1363514, -25'd4834275, -25'd991646, -25'd3718673, 25'd206593}, '{-25'd454505, -25'd3842629, 25'd4669001, -25'd1404832, -25'd3057576, -25'd1776699, 25'd909009, 25'd2520434, 25'd2561753}, '{-25'd661097, 25'd2355160, -25'd495823, 25'd3759992, -25'd4421089, -25'd2685709, 25'd2974939, -25'd1776699, 25'd3057576}, '{-25'd165274, 25'd3470762, -25'd123956, -25'd1363514, -25'd4462408, 25'd2933620, -25'd1032965, -25'd2479116, -25'd3512080}, '{25'd2479116, -25'd3594718, -25'd4710320, -25'd4338452, 25'd1528788, 25'd826372, 25'd1198239, 25'd1735381, 25'd1322195}}, '{'{-25'd2768346, -25'd3222850, 25'd4007903, -25'd3553399, -25'd3925266, 25'd2892301, -25'd1941974, -25'd3057576, 25'd2479116}, '{25'd2727027, 25'd2603071, -25'd1818018, 25'd4669001, 25'd2024611, -25'd4131859, 25'd2809664, -25'd247912, 25'd3842629}, '{-25'd1859337, -25'd4090541, 25'd3057576, 25'd1570107, 25'd5164824, -25'd3264169, 25'd1570107, -25'd1322195, -25'd661097}, '{-25'd2561753, -25'd4297134, 25'd4173178, 25'd1322195, 25'd2148567, 25'd4710320, 25'd2479116, 25'd2231204, 25'd3759992}, '{-25'd247912, 25'd4958231, 25'd3842629, -25'd4297134, 25'd2603071, 25'd2685709, -25'd1280876, 25'd2892301, -25'd247912}, '{25'd247912, 25'd2231204, 25'd2974939, -25'd4586364, 25'd2189885, -25'd1032965, -25'd2437797, -25'd2024611, 25'd1900655}, '{25'd3636036, -25'd1156921, -25'd3470762, -25'd3057576, 25'd2644390, 25'd2727027, 25'd5082187, 25'd1941974, 25'd3883948}, '{-25'd3305487, -25'd4421089, 25'd3346806, 25'd785053, 25'd743735, 25'd2644390, 25'd82637, 25'd1239558, -25'd950328}, '{25'd2561753, 25'd3016257, 25'd1611425, 25'd247912, -25'd3718673, -25'd454505, 25'd2561753, -25'd1528788, 25'd3925266}}},
    '{'{'{-25'd1368092, -25'd1809413, -25'd882640, 25'd3221637, -25'd1191564, 25'd485452, 25'd2294865, -25'd1015036, -25'd3707089}, '{25'd2294865, -25'd3530561, 25'd3309901, -25'd4104277, -25'd3045109, -25'd4898654, -25'd4280805, -25'd308924, -25'd573716}, '{25'd1500488, -25'd661980, 25'd2471393, -25'd2074205, 25'd4060145, 25'd3618825, 25'd485452, 25'd1456356, -25'd3662957}, '{-25'd4545597, -25'd132396, 25'd3662957, -25'd3486429, -25'd4457333, 25'd4413201, -25'd4854522, 25'd485452, 25'd2030073}, '{-25'd3662957, 25'd397188, 25'd4060145, -25'd3662957, -25'd2383129, -25'd44132, -25'd3133373, -25'd5119314, 25'd1853545}, '{-25'd529584, 25'd2692053, -25'd3662957, -25'd4192541, -25'd3839485, 25'd3618825, -25'd1544621, 25'd882640, -25'd3486429}, '{-25'd3000977, 25'd2206601, -25'd3751221, -25'd3309901, 25'd2956845, 25'd2824449, 25'd2030073, 25'd4413201, 25'd2868581}, '{-25'd1500488, 25'd1500488, 25'd2647921, -25'd1897677, 25'd3883617, 25'd3662957, 25'd4324937, -25'd4236673, -25'd88264}, '{25'd2824449, -25'd4236673, 25'd3000977, 25'd1191564, 25'd1191564, -25'd5119314, 25'd4104277, -25'd3133373, 25'd2824449}}, '{'{-25'd3354033, 25'd926772, -25'd4016013, 25'd1279828, 25'd1588753, -25'd4148409, 25'd3618825, 25'd4104277, 25'd1588753}, '{25'd2338997, -25'd4192541, 25'd1677017, -25'd441320, 25'd2118337, -25'd5031050, -25'd4501465, 25'd706112, -25'd2868581}, '{-25'd2162469, -25'd4722126, -25'd4457333, 25'd3398165, 25'd441320, -25'd2868581, -25'd1721149, -25'd485452, 25'd3398165}, '{25'd3177505, -25'd5163446, -25'd4722126, -25'd2383129, 25'd1279828, -25'd1941809, -25'd4589730, -25'd3045109, 25'd750244}, '{-25'd4545597, -25'd1059168, -25'd3530561, -25'd4854522, 25'd1677017, 25'd2956845, 25'd1765281, -25'd4192541, 25'd2118337}, '{-25'd1279828, -25'd794376, -25'd750244, -25'd2206601, -25'd794376, -25'd441320, 25'd2383129, -25'd750244, -25'd4413201}, '{25'd2515525, 25'd4236673, -25'd3751221, 25'd4501465, 25'd3354033, 25'd3751221, 25'd2515525, -25'd1368092, -25'd1765281}, '{25'd2338997, 25'd2868581, 25'd3221637, 25'd3574693, 25'd3883617, -25'd2427261, 25'd3971881, -25'd926772, 25'd2736185}, '{-25'd220660, -25'd2162469, 25'd2515525, 25'd661980, 25'd4457333, -25'd2383129, -25'd4810390, 25'd3618825, -25'd1323960}}, '{'{-25'd308924, -25'd44132, -25'd4854522, -25'd5031050, 25'd4501465, 25'd2603789, -25'd3221637, -25'd44132, 25'd4457333}, '{-25'd5604766, -25'd5604766, -25'd5648898, 25'd3574693, 25'd1456356, 25'd3751221, -25'd4854522, 25'd2250733, -25'd4986918}, '{-25'd3354033, 25'd308924, 25'd1191564, 25'd882640, 25'd3398165, 25'd4501465, 25'd3751221, -25'd3265769, -25'd4148409}, '{25'd3354033, -25'd1853545, -25'd3839485, 25'd3486429, 25'd3707089, 25'd1103300, 25'd4016013, 25'd4501465, 25'd3574693}, '{-25'd3133373, 25'd1235696, 25'd176528, 25'd661980, -25'd4898654, 25'd2515525, -25'd4236673, 25'd4457333, 25'd970904}, '{25'd838508, -25'd617848, 25'd3133373, 25'd2956845, 25'd2338997, 25'd970904, 25'd2074205, 25'd4589730, 25'd2427261}, '{-25'd3045109, 25'd3751221, 25'd264792, 25'd3971881, -25'd3971881, 25'd1412224, -25'd2383129, -25'd4810390, -25'd1853545}, '{25'd2030073, -25'd1632885, -25'd2383129, 25'd2780317, -25'd3839485, -25'd3662957, 25'd4324937, 25'd1191564, -25'd4589730}, '{-25'd176528, 25'd661980, -25'd882640, 25'd44132, 25'd1985941, -25'd1191564, -25'd3177505, -25'd794376, -25'd2824449}}},
    '{'{'{25'd376184, 25'd2006315, 25'd4388814, -25'd4221621, 25'd3260262, -25'd4263419, 25'd1880920, 25'd3720042, 25'd4723199}, '{25'd4054428, -25'd4305217, 25'd1003157, 25'd835965, -25'd4388814, 25'd2758683, 25'd3218463, 25'd1546534, 25'd1044956}, '{25'd4388814, 25'd3511051, -25'd752368, -25'd3720042, -25'd4514208, 25'd3302060, 25'd877763, 25'd752368, -25'd2257104}, '{25'd585175, -25'd83596, -25'd501579, -25'd1546534, 25'd1504736, -25'd1671929, -25'd3260262, -25'd4138024, 25'd3636446}, '{-25'd1671929, -25'd2382499, 25'd334386, -25'd961359, -25'd835965, -25'd1337543, -25'd3260262, -25'd292588, 25'd961359}, '{-25'd2633288, 25'd835965, -25'd41798, 25'd794166, 25'd2215306, -25'd2424297, -25'd1086754, 25'd2675086, -25'd1253947}, '{-25'd417982, -25'd4764998, 25'd417982, 25'd2466095, -25'd3511051, 25'd3093069, -25'd2006315, 25'd3845437, 25'd3051270}, '{25'd208991, -25'd2298902, 25'd3594647, 25'd2089911, 25'd2591490, 25'd1839122, -25'd3218463, 25'd167193, -25'd4932191}, '{25'd2925876, 25'd3427454, 25'd835965, 25'd2884078, -25'd3970831, 25'd459780, 25'd1253947, 25'd4639603, -25'd376184}}, '{'{25'd1630131, -25'd1797324, 25'd1713727, -25'd501579, -25'd3594647, 25'd208991, -25'd1003157, -25'd3134867, 25'd3260262}, '{-25'd2842279, -25'd1253947, -25'd3093069, -25'd1003157, -25'd2340701, 25'd501579, 25'd877763, 25'd1170350, 25'd3218463}, '{-25'd2507894, 25'd1253947, -25'd4639603, -25'd2048113, -25'd1922718, 25'd1504736, -25'd2257104, 25'd2549692, -25'd961359}, '{-25'd5266576, -25'd125395, 25'd1671929, 25'd835965, 25'd4096226, -25'd1170350, -25'd459780, 25'd0, 25'd4054428}, '{25'd4472410, -25'd877763, -25'd1086754, -25'd2257104, 25'd3970831, -25'd5308375, 25'd3093069, 25'd961359, -25'd1630131}, '{-25'd4597805, -25'd2800481, -25'd334386, 25'd2967674, -25'd626973, 25'd2131709, -25'd1462938, 25'd1253947, -25'd1086754}, '{25'd3761840, 25'd585175, 25'd3636446, -25'd2842279, -25'd5350173, 25'd3302060, 25'd1964517, -25'd3469253, -25'd877763}, '{25'd961359, 25'd2048113, 25'd208991, -25'd2298902, 25'd3218463, 25'd543377, -25'd1504736, 25'd2758683, -25'd961359}, '{-25'd459780, -25'd501579, 25'd2298902, -25'd2925876, -25'd208991, 25'd3093069, -25'd1797324, 25'd4054428, 25'd1003157}}, '{'{-25'd4764998, -25'd3887235, 25'd2800481, -25'd2591490, 25'd4347015, 25'd3845437, -25'd1379341, -25'd1630131, -25'd2131709}, '{-25'd1839122, -25'd3051270, 25'd2089911, -25'd2131709, -25'd4514208, 25'd585175, -25'd4138024, 25'd4973989, 25'd626973}, '{25'd4430612, 25'd1379341, -25'd752368, -25'd5057585, 25'd3385656, -25'd1044956, 25'd208991, -25'd1588333, -25'd501579}, '{-25'd459780, 25'd4514208, -25'd3552849, 25'd1504736, 25'd4054428, 25'd1170350, -25'd585175, 25'd2675086, -25'd3051270}, '{25'd4179823, 25'd3929033, -25'd376184, 25'd543377, 25'd1504736, 25'd2591490, 25'd4347015, -25'd167193, 25'd2048113}, '{25'd1964517, 25'd3552849, 25'd3970831, -25'd2466095, 25'd919561, -25'd3302060, 25'd1295745, 25'd3218463, 25'd710570}, '{-25'd2298902, 25'd2800481, 25'd1003157, -25'd2925876, -25'd710570, -25'd877763, 25'd4597805, -25'd752368, -25'd2048113}, '{25'd2758683, -25'd3176665, -25'd961359, 25'd208991, 25'd1630131, 25'd2925876, 25'd961359, -25'd4848594, 25'd668772}, '{-25'd4681401, 25'd2967674, 25'd3176665, 25'd3051270, 25'd4890392, 25'd4514208, -25'd125395, 25'd3009472, 25'd4179823}}},
    '{'{'{-25'd2064474, -25'd2223280, 25'd3890740, -25'd794029, -25'd4605366, 25'd2739399, -25'd3890740, 25'd4208352, 25'd4565664}, '{-25'd4446560, -25'd3454024, -25'd2183579, 25'd3136413, 25'd317611, 25'd1985072, 25'd754327, 25'd714626, 25'd4605366}, '{-25'd1985072, -25'd4446560, -25'd1032237, -25'd3652532, 25'd2461489, 25'd3692233, -25'd1191043, 25'd635223, 25'd317611}, '{-25'd3533427, -25'd4883276, -25'd158806, 25'd2977607, -25'd2024773, 25'd1349849, 25'd4009844, -25'd3096712, 25'd1111640}, '{25'd4049546, -25'd3454024, 25'd1310147, 25'd4287754, 25'd2818802, -25'd3612830, -25'd3334920, 25'd4406859, 25'd1468953}, '{25'd3334920, 25'd635223, -25'd3890740, 25'd5042082, -25'd952834, 25'd4287754, 25'd3493726, -25'd2977607, 25'd4287754}, '{-25'd3652532, 25'd4565664, 25'd1548356, 25'd2302683, -25'd277910, 25'd3731934, 25'd39701, -25'd119104, -25'd4724470}, '{-25'd3295219, -25'd4208352, 25'd3255517, 25'd4367157, 25'd1985072, -25'd1468953, 25'd2064474, -25'd3493726, 25'd4486262}, '{-25'd397014, -25'd4168650, -25'd3295219, -25'd4486262, 25'd2064474, -25'd1389550, -25'd3771636, -25'd1429251, 25'd2739399}}, '{'{25'd2421787, -25'd2580593, 25'd3851039, 25'd3612830, -25'd4406859, -25'd2104176, -25'd4843575, -25'd1508654, 25'd1826266}, '{25'd3533427, 25'd4605366, 25'd2620294, -25'd1349849, -25'd1826266, 25'd3057010, 25'd2262982, 25'd2183579, -25'd2183579}, '{25'd4843575, -25'd158806, 25'd1707162, -25'd3295219, 25'd476417, -25'd158806, -25'd3454024, -25'd476417, -25'd3573129}, '{-25'd833730, -25'd4645067, -25'd2223280, 25'd1786564, 25'd436716, 25'd1627759, 25'd1389550, 25'd3533427, -25'd3414323}, '{-25'd3652532, -25'd1349849, -25'd1786564, -25'd1826266, 25'd952834, 25'd2302683, 25'd277910, 25'd1865967, 25'd754327}, '{25'd2540892, -25'd1111640, 25'd317611, 25'd3731934, 25'd4565664, 25'd2382086, -25'd1468953, -25'd4803873, -25'd635223}, '{25'd3493726, -25'd595521, 25'd2977607, 25'd4009844, 25'd4605366, 25'd2104176, 25'd4208352, 25'd754327, 25'd1151341}, '{-25'd1270446, 25'd4525963, 25'd2382086, 25'd3096712, -25'd2699697, -25'd952834, -25'd1349849, -25'd2977607, -25'd2143877}, '{-25'd2898204, 25'd2183579, -25'd1627759, 25'd2104176, -25'd1588057, -25'd4367157, -25'd833730, 25'd1746863, 25'd4168650}}, '{'{-25'd952834, -25'd4248053, 25'd833730, -25'd1230744, 25'd1389550, -25'd119104, -25'd1191043, 25'd119104, 25'd4446560}, '{-25'd4446560, -25'd4724470, 25'd2937906, 25'd1389550, -25'd4446560, 25'd476417, -25'd4922977, 25'd1310147, 25'd4208352}, '{25'd913133, -25'd2223280, 25'd2937906, 25'd1071939, 25'd397014, -25'd317611, -25'd39701, -25'd635223, -25'd4565664}, '{25'd436716, 25'd1111640, -25'd1071939, 25'd2382086, -25'd3295219, -25'd3414323, -25'd1032237, 25'd3255517, -25'd2620294}, '{25'd754327, 25'd1627759, -25'd2183579, 25'd1349849, 25'd158806, 25'd1627759, 25'd317611, 25'd4168650, 25'd3573129}, '{25'd3811337, -25'd1270446, -25'd3017309, 25'd3295219, 25'd833730, -25'd2461489, -25'd2461489, 25'd1071939, 25'd1349849}, '{-25'd1151341, -25'd3255517, 25'd1032237, 25'd2262982, 25'd913133, -25'd79403, -25'd1667460, -25'd2342384, -25'd595521}, '{-25'd674924, 25'd3851039, 25'd4803873, 25'd2501190, 25'd3612830, 25'd4208352, -25'd2461489, 25'd2540892, -25'd4009844}, '{-25'd3652532, -25'd1230744, -25'd2858503, 25'd3057010, -25'd4962679, -25'd3454024, -25'd3295219, 25'd2104176, 25'd1508654}}},
    '{'{'{-25'd2677841, 25'd167365, 25'd2217587, -25'd2552318, 25'd209206, -25'd669460, -25'd1966540, 25'd4769905, -25'd3054413}, '{25'd3138095, 25'd1548127, 25'd2761524, 25'd2384953, -25'd585778, 25'd585778, 25'd2677841, 25'd2092064, 25'd920508}, '{-25'd83683, 25'd2636000, 25'd292889, -25'd3472826, 25'd2594159, 25'd1004191, 25'd2175746, -25'd2510476, 25'd4937270}, '{-25'd2552318, 25'd4184127, 25'd794984, -25'd1506286, -25'd418413, -25'd1589968, -25'd1548127, 25'd1631810, -25'd920508}, '{25'd1171556, -25'd2887048, -25'd3096254, 25'd1882857, 25'd5104635, -25'd2887048, 25'd1380762, -25'd3598349, 25'd4602540}, '{-25'd3807556, 25'd1673651, 25'd2259429, 25'd5313842, 25'd4351492, 25'd2384953, 25'd4184127, -25'd3974921, 25'd3598349}, '{25'd2175746, -25'd2887048, -25'd2133905, -25'd3221778, 25'd251048, -25'd125524, -25'd1882857, -25'd3807556, -25'd2426794}, '{25'd3430984, 25'd2426794, 25'd3179937, 25'd0, 25'd585778, -25'd3974921, 25'd2677841, 25'd4895429, -25'd4435175}, '{25'd3640191, 25'd3263619, 25'd4435175, 25'd3974921, -25'd4100445, 25'd1464445, -25'd962349, 25'd2217587, 25'd4979111}}, '{'{25'd836825, 25'd1841016, -25'd794984, -25'd41841, 25'd334730, -25'd3054413, 25'd1631810, 25'd3556508, 25'd2510476}, '{-25'd1589968, 25'd2552318, -25'd3598349, -25'd3933080, -25'd4518857, 25'd502095, 25'd2008381, 25'd2050222, -25'd4728064}, '{-25'd2928889, 25'd4393334, 25'd3096254, -25'd2970730, 25'd2384953, -25'd167365, 25'd4184127, -25'd3430984, 25'd1422603}, '{25'd3138095, -25'd2636000, -25'd3472826, 25'd1129714, 25'd5020953, -25'd376571, 25'd3430984, 25'd3807556, -25'd1841016}, '{-25'd3221778, 25'd4811746, 25'd3305461, 25'd2677841, 25'd4602540, 25'd2217587, 25'd292889, -25'd3012572, -25'd3682032}, '{-25'd4309651, 25'd3682032, 25'd1004191, 25'd2719683, -25'd4225969, 25'd2928889, -25'd2761524, -25'd209206, 25'd2677841}, '{25'd4644381, 25'd2008381, -25'd1046032, -25'd4435175, -25'd2594159, -25'd3221778, 25'd1129714, -25'd3974921, -25'd3263619}, '{-25'd2133905, 25'd2510476, 25'd920508, 25'd418413, 25'd2259429, 25'd3598349, -25'd2343111, -25'd1841016, 25'd1631810}, '{25'd83683, 25'd1966540, -25'd4811746, -25'd3556508, -25'd251048, -25'd1631810, -25'd794984, 25'd1548127, -25'd460254}}, '{'{25'd3723873, 25'd3472826, -25'd3472826, -25'd4351492, -25'd1464445, 25'd2217587, 25'd1548127, -25'd3347302, 25'd3891238}, '{-25'd1882857, 25'd4309651, 25'd836825, 25'd4686223, -25'd3640191, -25'd2133905, -25'd2677841, -25'd836825, -25'd3221778}, '{-25'd3807556, -25'd1882857, 25'd41841, -25'd418413, 25'd3974921, 25'd3389143, -25'd2719683, -25'd3138095, -25'd4728064}, '{-25'd2636000, -25'd125524, 25'd3347302, 25'd1882857, 25'd2803365, 25'd5020953, -25'd1715492, -25'd167365, 25'd2092064}, '{25'd1213397, 25'd4309651, 25'd2636000, -25'd209206, 25'd4560699, -25'd4184127, 25'd3012572, 25'd1548127, -25'd4225969}, '{25'd669460, 25'd4100445, 25'd1422603, 25'd125524, -25'd2552318, -25'd1589968, 25'd209206, -25'd1213397, -25'd502095}, '{25'd251048, 25'd1506286, -25'd1757333, -25'd3221778, -25'd2970730, 25'd1715492, 25'd167365, -25'd1255238, 25'd3179937}, '{25'd4058603, -25'd4100445, -25'd3263619, 25'd3179937, -25'd3933080, 25'd585778, -25'd3598349, 25'd4769905, -25'd3389143}, '{25'd3347302, -25'd4435175, 25'd4016762, 25'd3054413, 25'd1506286, 25'd460254, 25'd83683, -25'd4225969, -25'd1422603}}},
    '{'{'{-25'd3075811, 25'd958040, -25'd3126234, -25'd857193, 25'd4487659, -25'd4840621, 25'd1361425, 25'd1411848, 25'd554654}, '{25'd3580042, -25'd1411848, -25'd3277504, 25'd605078, -25'd3327927, -25'd907616, 25'd201693, -25'd2117772, 25'd3630465}, '{-25'd4235543, -25'd1109309, 25'd3378350, -25'd1563117, 25'd806770, 25'd2369887, 25'd1260578, 25'd958040, -25'd4185120}, '{-25'd4235543, 25'd453808, -25'd1966502, 25'd5697814, 25'd6403738, 25'd4437236, 25'd4134697, -25'd806770, -25'd1966502}, '{-25'd605078, 25'd2218618, 25'd2117772, 25'd6403738, 25'd4538082, 25'd806770, -25'd1311001, 25'd302539, -25'd5143159}, '{-25'd4084274, -25'd1109309, -25'd504231, 25'd1058886, 25'd554654, -25'd6454161, 25'd0, 25'd1815233, -25'd4991890}, '{-25'd1663963, 25'd1613540, 25'd3680889, -25'd3781735, -25'd2117772, -25'd6050776, -25'd2016925, -25'd2672426, 25'd2117772}, '{-25'd1815233, -25'd3731312, -25'd2672426, 25'd2420310, -25'd3983427, -25'd2672426, -25'd2571580, 25'd1058886, 25'd3479196}, '{-25'd907616, -25'd151269, -25'd100846, 25'd2218618, -25'd2319464, -25'd50423, -25'd2571580, 25'd2874119, 25'd2016925}}, '{'{25'd3479196, 25'd3882581, -25'd3227080, -25'd1210155, -25'd403385, 25'd1008463, 25'd1714386, -25'd1058886, 25'd958040}, '{-25'd3529619, 25'd5445698, -25'd1663963, -25'd2016925, -25'd1462271, -25'd1966502, 25'd4285966, -25'd5092736, 25'd1210155}, '{25'd2470733, 25'd151269, -25'd1109309, 25'd3025388, 25'd3781735, -25'd1008463, -25'd1865656, 25'd151269, -25'd3126234}, '{-25'd958040, -25'd3580042, 25'd3731312, 25'd0, 25'd3630465, -25'd3126234, -25'd806770, -25'd5042313, 25'd705924}, '{-25'd50423, -25'd705924, -25'd1008463, 25'd4033851, 25'd4336389, 25'd5748237, 25'd1411848, -25'd554654, -25'd3075811}, '{-25'd2420310, 25'd3378350, -25'd2672426, 25'd2924542, -25'd1058886, -25'd2672426, -25'd1563117, 25'd2319464, -25'd5042313}, '{-25'd5294429, 25'd504231, -25'd1462271, -25'd3781735, -25'd252116, -25'd5344852, 25'd907616, -25'd3277504, -25'd705924}, '{25'd252116, -25'd1058886, 25'd302539, -25'd2974965, -25'd3781735, -25'd857193, -25'd5042313, -25'd1058886, 25'd3680889}, '{-25'd2168195, -25'd2924542, 25'd4689351, -25'd4538082, 25'd504231, 25'd3227080, -25'd2823695, 25'd2773272, 25'd4285966}}, '{'{25'd3983427, 25'd2521157, -25'd100846, 25'd504231, -25'd554654, -25'd6050776, -25'd6252468, -25'd5949930, -25'd4185120}, '{-25'd3378350, -25'd756347, -25'd605078, 25'd3731312, 25'd2168195, -25'd1411848, -25'd3832158, -25'd3731312, 25'd0}, '{-25'd1916079, 25'd50423, 25'd1058886, -25'd2672426, 25'd5143159, -25'd3580042, 25'd2016925, -25'd2722849, 25'd2924542}, '{-25'd554654, -25'd4739774, 25'd3580042, 25'd958040, 25'd3781735, 25'd655501, 25'd1663963, -25'd3428773, -25'd1260578}, '{-25'd4386812, -25'd806770, 25'd3277504, 25'd2722849, 25'd5849083, -25'd857193, -25'd3075811, -25'd3277504, 25'd3428773}, '{25'd100846, 25'd1512694, -25'd4991890, 25'd3933004, -25'd1411848, -25'd1311001, -25'd2016925, 25'd4689351, -25'd4739774}, '{-25'd5496121, 25'd2622003, -25'd2823695, 25'd1159732, 25'd2672426, -25'd201693, 25'd1058886, 25'd302539, 25'd352962}, '{-25'd3479196, -25'd1764810, -25'd3479196, -25'd1210155, 25'd1865656, 25'd3680889, -25'd3781735, 25'd3882581, 25'd1008463}, '{25'd3378350, 25'd2874119, -25'd1411848, -25'd3731312, 25'd1966502, -25'd5849083, -25'd806770, -25'd252116, 25'd4891044}}},
    '{'{'{25'd556312, -25'd3295080, -25'd641899, -25'd4750051, -25'd2225249, 25'd3894186, -25'd2824355, -25'd1626144, 25'd385139}, '{25'd2695975, -25'd2396422, 25'd3551840, -25'd1626144, 25'd4150945, -25'd2952734, -25'd2182456, -25'd4536085, -25'd2952734}, '{25'd1326591, -25'd3680220, -25'd3808599, 25'd4193739, 25'd3423460, 25'd1155418, 25'd2054076, -25'd4964017, 25'd3380667}, '{25'd1711730, 25'd3123907, 25'd2182456, 25'd2396422, 25'd2995528, -25'd2225249, 25'd1412177, -25'd85587, 25'd3637426}, '{-25'd4364912, -25'd3680220, 25'd2995528, -25'd5135190, -25'd4792844, -25'd2995528, 25'd2867148, -25'd4964017, 25'd3423460}, '{25'd1968490, -25'd641899, -25'd5177983, -25'd1283798, -25'd1369384, 25'd2268042, 25'd3209494, -25'd2011283, -25'd4065359}, '{-25'd727485, -25'd2524802, 25'd3894186, 25'd4407705, -25'd2909941, 25'd1027038, -25'd2781561, 25'd3894186, -25'd1412177}, '{-25'd1069831, -25'd470726, 25'd941452, 25'd1155418, 25'd2182456, -25'd2995528, -25'd2439215, 25'd684692, 25'd3295080}, '{25'd85587, -25'd1840110, 25'd3380667, 25'd171173, -25'd3123907, 25'd4065359, -25'd3209494, -25'd3123907, -25'd4878431}}, '{'{-25'd5349156, -25'd3209494, -25'd984245, 25'd2439215, 25'd1241004, 25'd4150945, 25'd2054076, 25'd2482009, 25'd2396422}, '{25'd1711730, 25'd0, -25'd4493291, -25'd2738768, -25'd770279, 25'd4150945, -25'd1668937, 25'd855865, -25'd1369384}, '{-25'd3765806, -25'd684692, 25'd3808599, -25'd2268042, 25'd42793, 25'd1241004, 25'd1412177, 25'd898658, -25'd2738768}, '{-25'd256760, -25'd556312, 25'd3637426, 25'd3594633, -25'd1925696, -25'd4108152, 25'd2396422, -25'd3979772, 25'd1968490}, '{25'd2011283, -25'd1797317, -25'd1454971, -25'd4108152, -25'd1711730, -25'd684692, -25'd3252287, 25'd4621671, 25'd3081114}, '{25'd941452, 25'd2909941, 25'd1711730, -25'd2524802, 25'd2268042, 25'd1754523, -25'd2738768, -25'd4279325, 25'd1412177}, '{-25'd1968490, 25'd470726, 25'd4279325, -25'd1711730, -25'd1155418, -25'd4065359, 25'd1112625, -25'd5135190, -25'd4621671}, '{25'd941452, 25'd641899, -25'd2909941, -25'd3123907, 25'd1925696, 25'd3637426, 25'd4407705, -25'd213966, -25'd4578878}, '{25'd1711730, -25'd1583350, 25'd2396422, 25'd2653182, -25'd2054076, -25'd3637426, 25'd3337874, -25'd4022566, 25'd1668937}}, '{'{25'd1925696, -25'd5391950, -25'd3081114, 25'd2653182, 25'd2610388, -25'd1840110, -25'd813072, -25'd4493291, -25'd2738768}, '{-25'd5477536, -25'd1968490, 25'd1583350, -25'd2225249, -25'd5220777, -25'd5135190, -25'd4921224, 25'd1583350, 25'd4108152}, '{25'd2054076, -25'd5049604, -25'd4236532, 25'd3509047, -25'd2995528, -25'd2567595, -25'd4279325, 25'd941452, -25'd3081114}, '{25'd1882903, -25'd641899, 25'd4493291, -25'd2268042, -25'd3509047, 25'd4621671, 25'd2695975, -25'd1198211, 25'd3551840}, '{-25'd2096869, -25'd984245, -25'd256760, -25'd3723013, 25'd1369384, 25'd770279, 25'd556312, 25'd4878431, 25'd0}, '{25'd727485, 25'd3551840, 25'd3166701, 25'd299553, -25'd3123907, 25'd4022566, -25'd299553, 25'd213966, 25'd1668937}, '{-25'd1668937, 25'd4878431, -25'd1283798, 25'd2653182, 25'd2011283, -25'd3808599, -25'd1797317, -25'd2054076, 25'd2867148}, '{-25'd2225249, -25'd470726, -25'd2653182, 25'd3252287, 25'd4493291, 25'd4236532, 25'd1198211, -25'd470726, 25'd2867148}, '{25'd599106, 25'd3081114, 25'd4707258, -25'd2482009, 25'd4578878, 25'd3466253, 25'd2182456, 25'd4707258, 25'd2995528}}},
    '{'{'{-25'd921008, 25'd2930479, 25'd2846751, -25'd3767758, -25'd3516574, -25'd1465239, -25'd1716423, 25'd418640, -25'd2260655}, '{25'd1967607, 25'd502368, 25'd2218791, 25'd3056071, -25'd1381511, -25'd5358590, -25'd418640, 25'd962872, 25'd334912}, '{25'd2804887, 25'd1088464, -25'd4102670, -25'd4018942, 25'd376776, -25'd879144, -25'd2051335, -25'd3809622, 25'd418640}, '{-25'd3307254, 25'd2302519, -25'd4228262, -25'd3935214, -25'd1255919, 25'd2679295, 25'd921008, -25'd2428111, 25'd921008}, '{-25'd4772494, 25'd293048, 25'd5107406, 25'd2553703, 25'd544232, 25'd2428111, 25'd502368, 25'd1465239, 25'd837280}, '{-25'd3390982, 25'd4814358, -25'd1507103, 25'd2846751, 25'd3139799, -25'd2595567, 25'd460504, -25'd5358590, -25'd4939950}, '{25'd1339647, -25'd2135063, 25'd2972343, 25'd3390982, -25'd3600302, -25'd5358590, -25'd1590831, -25'd5358590, 25'd3432846}, '{25'd1842015, -25'd1590831, 25'd1423375, 25'd251184, -25'd5149270, -25'd4521310, -25'd837280, -25'd837280, 25'd460504}, '{-25'd1339647, 25'd251184, 25'd2260655, 25'd627960, -25'd2595567, -25'd5274862, -25'd2637431, 25'd753552, 25'd4437582}}, '{'{-25'd4688766, -25'd1465239, 25'd4898086, 25'd2511839, -25'd4186398, -25'd502368, 25'd2804887, 25'd1674559, -25'd1507103}, '{25'd0, -25'd1842015, 25'd3307254, 25'd2888615, 25'd1046600, 25'd3181663, -25'd5316726, 25'd209320, 25'd502368}, '{-25'd2302519, -25'd1046600, 25'd4939950, 25'd3977078, 25'd3474710, -25'd1758287, -25'd5358590, -25'd4395718, -25'd4353854}, '{25'd4563174, -25'd1339647, -25'd3181663, 25'd2595567, 25'd4856222, -25'd4437582, 25'd2469975, 25'd2386247, 25'd2176927}, '{25'd4939950, 25'd3935214, 25'd1339647, 25'd5316726, -25'd2846751, 25'd3181663, -25'd5358590, -25'd5191134, 25'd4772494}, '{25'd4437582, 25'd2679295, -25'd167456, -25'd209320, 25'd1088464, -25'd2093199, 25'd1883879, -25'd4144534, -25'd209320}, '{-25'd2386247, -25'd1465239, -25'd3390982, 25'd1716423, -25'd3181663, -25'd2972343, -25'd4856222, -25'd3977078, 25'd5316726}, '{-25'd3684030, -25'd4018942, -25'd1381511, 25'd2721159, -25'd3977078, -25'd2093199, -25'd2595567, 25'd1088464, 25'd5316726}, '{-25'd2135063, -25'd3893350, -25'd1842015, 25'd586096, -25'd4060806, -25'd4228262, -25'd1130327, 25'd4772494, 25'd5316726}}, '{'{25'd2428111, 25'd4688766, -25'd4437582, -25'd1548967, -25'd251184, -25'd1925743, -25'd1172191, -25'd753552, 25'd1967607}, '{-25'd2386247, 25'd4688766, -25'd1967607, 25'd4479446, -25'd3558438, 25'd3097935, -25'd1046600, 25'd3390982, -25'd586096}, '{25'd669824, -25'd334912, 25'd2637431, 25'd627960, 25'd125592, -25'd4521310, -25'd5107406, 25'd3684030, -25'd3307254}, '{-25'd83728, 25'd2930479, 25'd2972343, 25'd5316726, -25'd2218791, 25'd2093199, -25'd4186398, 25'd3432846, -25'd5107406}, '{-25'd2344383, -25'd293048, 25'd3809622, -25'd460504, -25'd1674559, -25'd3139799, -25'd4479446, 25'd2846751, -25'd4395718}, '{25'd753552, -25'd3014207, 25'd5149270, 25'd4688766, 25'd2428111, 25'd3223527, -25'd1088464, -25'd544232, 25'd5274862}, '{-25'd1800151, -25'd1214055, 25'd2763023, 25'd2511839, -25'd4605038, 25'd3181663, 25'd3851486, -25'd4270126, 25'd2093199}, '{25'd2721159, -25'd2721159, 25'd3642166, -25'd2637431, 25'd837280, -25'd1214055, -25'd209320, 25'd4898086, 25'd2846751}, '{25'd3014207, 25'd3014207, 25'd3684030, 25'd1297783, 25'd3307254, 25'd2218791, -25'd1925743, 25'd5316726, 25'd4730630}}},
    '{'{'{25'd760177, 25'd760177, -25'd1296773, -25'd2817127, 25'd3443156, -25'd1162624, -25'd4203333, 25'd2772411, -25'd2414681}, '{25'd268298, 25'd2369964, 25'd2146383, -25'd3711454, 25'd178865, -25'd2280532, 25'd536596, 25'd2280532, 25'd1565071}, '{-25'd2414681, 25'd4516347, 25'd2548830, 25'd804894, -25'd1341489, -25'd4471631, 25'd3622021, 25'd1162624, 25'd3264291}, '{-25'd3979752, -25'd3890319, -25'd1609787, -25'd2191099, 25'd1788652, 25'd5276524, -25'd1565071, 25'd2056950, -25'd2414681}, '{-25'd849610, -25'd983759, 25'd4963510, 25'd4292766, -25'd760177, 25'd1609787, 25'd3040709, 25'd4739929, 25'd536596}, '{25'd2682979, 25'd4203333, 25'd4024468, -25'd3130142, -25'd2951276, -25'd4561064, 25'd2772411, 25'd4024468, -25'd4248049}, '{-25'd5500106, -25'd313014, 25'd2280532, -25'd3666737, 25'd1609787, -25'd894326, -25'd3622021, 25'd2414681, -25'd1430922}, '{-25'd4784645, -25'd3935035, 25'd2459397, -25'd3935035, -25'd939042, -25'd5723688, -25'd1520355, -25'd4248049, 25'd0}, '{-25'd3040709, 25'd2951276, -25'd626028, -25'd4158617, 25'd3040709, -25'd3577305, -25'd5678971, -25'd44716, -25'd1117908}}, '{'{-25'd4874078, -25'd4471631, -25'd223582, 25'd1252057, -25'd2459397, -25'd2682979, 25'd2682979, -25'd3309007, -25'd4650496}, '{25'd1699220, 25'd3756170, -25'd849610, 25'd4292766, -25'd3577305, 25'd4874078, 25'd1967518, -25'd894326, -25'd89433}, '{-25'd2191099, 25'd1609787, -25'd2638262, -25'd4784645, -25'd3711454, -25'd357730, -25'd447163, -25'd1430922, 25'd3264291}, '{-25'd1743936, -25'd2995993, -25'd3309007, 25'd402447, 25'd2012234, 25'd4069184, 25'd357730, 25'd626028, -25'd3845603}, '{25'd2369964, -25'd1073191, 25'd4337482, 25'd5008227, -25'd3219574, -25'd4158617, -25'd1565071, 25'd3845603, 25'd1296773}, '{25'd402447, -25'd3040709, 25'd3622021, -25'd3040709, -25'd1520355, 25'd4069184, 25'd1520355, -25'd402447, -25'd2906560}, '{25'd134149, 25'd3577305, -25'd4158617, -25'd2995993, -25'd4650496, -25'd2593546, -25'd2235815, 25'd4337482, -25'd1028475}, '{-25'd4069184, -25'd3398440, -25'd2817127, -25'd2727695, 25'd715461, -25'd3577305, 25'd1609787, -25'd3219574, 25'd939042}, '{-25'd1565071, -25'd3085425, 25'd1162624, 25'd1296773, 25'd3353723, 25'd2682979, 25'd2682979, 25'd2817127, -25'd2548830}}, '{'{-25'd2995993, 25'd2056950, 25'd1699220, -25'd2414681, 25'd3040709, 25'd4158617, -25'd1162624, 25'd3577305, 25'd1609787}, '{-25'd760177, 25'd89433, -25'd44716, -25'd4337482, 25'd1967518, -25'd4248049, 25'd3443156, 25'd223582, -25'd3040709}, '{-25'd4918794, -25'd1654503, 25'd2861844, 25'd491879, -25'd1117908, 25'd4650496, -25'd357730, 25'd2280532, 25'd3487872}, '{25'd2682979, 25'd134149, -25'd2056950, 25'd3264291, -25'd2593546, -25'd3577305, -25'd44716, 25'd3890319, -25'd4471631}, '{25'd849610, -25'd3711454, -25'd1520355, -25'd1207340, 25'd894326, -25'd1833369, -25'd2817127, 25'd2012234, -25'd3711454}, '{-25'd1475638, -25'd5097659, -25'd1878085, -25'd4337482, 25'd2995993, 25'd626028, -25'd2995993, 25'd1341489, -25'd1788652}, '{25'd178865, 25'd89433, 25'd3487872, -25'd2861844, -25'd2593546, 25'd3622021, 25'd223582, 25'd89433, -25'd894326}, '{25'd1207340, -25'd4203333, 25'd1609787, 25'd4248049, 25'd313014, 25'd581312, 25'd4024468, 25'd5678971, 25'd4337482}, '{25'd3577305, -25'd2235815, -25'd3622021, 25'd1520355, -25'd2369964, 25'd3622021, 25'd2191099, -25'd3085425, -25'd2682979}}},
    '{'{'{25'd2020108, 25'd2772697, -25'd752589, -25'd4990855, -25'd4159046, -25'd4317485, -25'd4594755, -25'd3762946, -25'd2535037}, '{25'd1465568, 25'd2138938, -25'd3683726, -25'd2733087, 25'd118830, 25'd2099328, 25'd1901278, -25'd594149, 25'd4198656}, '{25'd2891527, -25'd4594755, -25'd2455817, 25'd2653867, -25'd2891527, -25'd1505178, 25'd2376597, 25'd158440, 25'd792199}, '{-25'd911029, 25'd4119436, 25'd3049967, -25'd3921386, 25'd1822058, 25'd1742838, 25'd3723336, -25'd4000606, 25'd990249}, '{25'd4713585, 25'd4198656, 25'd1227909, 25'd2693477, -25'd3723336, -25'd2535037, -25'd4673975, -25'd3406456, 25'd1663618}, '{25'd3683726, -25'd2416207, -25'd237660, -25'd1742838, 25'd316880, -25'd4357095, -25'd3248017, 25'd2535037, 25'd4159046}, '{25'd2614257, -25'd4634365, 25'd2059718, -25'd2931137, 25'd1307129, 25'd3525286, -25'd4673975, -25'd3842166, -25'd3485676}, '{-25'd2891527, -25'd4317485, -25'd4277875, -25'd1346739, 25'd2733087, 25'd3960996, -25'd3960996, -25'd1346739, -25'd2416207}, '{25'd2336988, 25'd2336988, 25'd831809, -25'd514929, 25'd2059718, 25'd1505178, -25'd1980498, -25'd2376597, 25'd2653867}}, '{'{-25'd316880, -25'd1742838, -25'd3604506, -25'd3446066, -25'd1069469, -25'd1703228, -25'd990249, -25'd3168797, -25'd1584398}, '{25'd3248017, -25'd3762946, -25'd911029, 25'd2614257, -25'd2178548, -25'd1425958, -25'd4436315, 25'd4238265, -25'd950639}, '{25'd435710, -25'd4634365, -25'd871419, -25'd3842166, -25'd2495427, 25'd237660, 25'd2297378, 25'd2257768, -25'd2772697}, '{-25'd990249, 25'd1703228, -25'd4119436, 25'd831809, -25'd3683726, 25'd1822058, -25'd39610, 25'd4713585, 25'd2218158}, '{-25'd2733087, 25'd79220, 25'd871419, 25'd1822058, 25'd2416207, -25'd3287626, 25'd39610, -25'd3960996, 25'd4396705}, '{-25'd39610, 25'd475319, 25'd3287626, -25'd2812307, 25'd3802556, 25'd3208407, -25'd2059718, 25'd118830, -25'd950639}, '{25'd277270, 25'd673369, 25'd3960996, -25'd1940888, 25'd1742838, -25'd4832415, 25'd79220, -25'd3723336, -25'd3644116}, '{25'd3366846, -25'd2812307, 25'd356490, -25'd831809, -25'd4951245, -25'd1980498, -25'd4832415, -25'd3168797, 25'd752589}, '{25'd1782448, -25'd554539, 25'd2495427, -25'd831809, -25'd2614257, 25'd4555145, -25'd118830, -25'd3525286, -25'd2891527}}, '{'{-25'd1822058, -25'd1703228, 25'd4198656, 25'd1584398, -25'd4832415, -25'd237660, -25'd3723336, -25'd1940888, 25'd1505178}, '{25'd2257768, 25'd4079826, 25'd594149, -25'd198050, -25'd4753195, 25'd1901278, 25'd3762946, -25'd4000606, -25'd1782448}, '{25'd4079826, -25'd2772697, 25'd1227909, -25'd3129187, 25'd2455817, 25'd2851917, 25'd2653867, 25'd3248017, -25'd792199}, '{25'd4634365, -25'd3406456, 25'd1109079, -25'd3683726, 25'd1544788, 25'd2138938, 25'd2812307, 25'd1425958, -25'd752589}, '{25'd2020108, -25'd2693477, 25'd1980498, -25'd2574647, 25'd514929, 25'd1663618, -25'd1782448, 25'd3525286, 25'd3208407}, '{-25'd1148689, 25'd3208407, 25'd911029, 25'd712979, -25'd4238265, -25'd1505178, -25'd2138938, -25'd237660, -25'd79220}, '{25'd2733087, 25'd633759, -25'd1069469, -25'd5070075, 25'd3644116, 25'd1307129, -25'd1624008, 25'd4792805, 25'd3683726}, '{-25'd4357095, -25'd2059718, 25'd1267519, -25'd4396705, -25'd2336988, -25'd4357095, -25'd2455817, 25'd1188299, -25'd1148689}, '{-25'd4951245, -25'd4911635, -25'd4713585, -25'd554539, 25'd3683726, 25'd3683726, 25'd158440, 25'd3049967, -25'd3960996}}},
    '{'{'{-25'd2175231, -25'd4350463, 25'd2835570, 25'd3068630, -25'd1903328, 25'd3962029, -25'd971085, -25'd4622367, -25'd3185160}, '{25'd1825641, -25'd427278, 25'd4233933, -25'd1709110, -25'd504964, 25'd4039716, 25'd4700054, -25'd4350463, 25'd3418221}, '{25'd2175231, 25'd2330605, -25'd971085, -25'd4117402, 25'd2952100, -25'd1592580, 25'd1165303, 25'd3923185, 25'd1942171}, '{-25'd621495, 25'd3457064, 25'd3651281, 25'd2835570, 25'd3340534, -25'd1553737, 25'd1165303, 25'd1048772, 25'd1126459}, '{25'd1903328, 25'd3340534, -25'd2641352, 25'd3495908, -25'd77687, -25'd2952100, 25'd3962029, -25'd4078559, 25'd4816584}, '{25'd4156246, -25'd2291762, -25'd738025, -25'd971085, 25'd4078559, -25'd2835570, 25'd3923185, 25'd2952100, -25'd4272776}, '{25'd1359520, 25'd271904, -25'd543808, 25'd1786797, 25'd4078559, 25'd194217, 25'd2874413, 25'd1514893, -25'd4505837}, '{25'd4233933, 25'd0, 25'd1087616, 25'd2447135, 25'd893399, -25'd4117402, 25'd2408292, 25'd4505837, 25'd3457064}, '{-25'd621495, -25'd2680196, -25'd2291762, 25'd1864484, -25'd1553737, -25'd2796726, -25'd3107473, -25'd2874413, 25'd4700054}}, '{'{25'd582651, 25'd776868, -25'd3146317, -25'd4544680, -25'd1631424, 25'd660338, -25'd3379377, 25'd3457064, 25'd2019858}, '{25'd2602509, 25'd2719039, 25'd3185160, 25'd1359520, -25'd1981014, 25'd3612438, -25'd2990943, 25'd2641352, -25'd543808}, '{-25'd271904, -25'd4195089, -25'd3379377, 25'd1087616, 25'd2175231, 25'd2874413, 25'd1009929, -25'd194217, 25'd1048772}, '{-25'd738025, -25'd3767812, 25'd2952100, -25'd466121, 25'd3806655, 25'd3379377, 25'd1242989, -25'd2369449, 25'd388434}, '{-25'd3651281, 25'd1437206, 25'd4777740, 25'd4894271, -25'd1126459, -25'd271904, -25'd3418221, -25'd3923185, 25'd1165303}, '{25'd621495, 25'd660338, 25'd971085, -25'd2641352, -25'd1165303, -25'd1009929, -25'd2719039, 25'd1592580, 25'd3612438}, '{25'd4428150, -25'd660338, -25'd427278, 25'd1747954, 25'd4894271, -25'd2136388, -25'd116530, 25'd3573594, 25'd1981014}, '{25'd2252918, 25'd2330605, 25'd2952100, 25'd776868, -25'd2136388, -25'd2136388, -25'd776868, 25'd2563666, 25'd1398363}, '{25'd1087616, 25'd4389306, -25'd2602509, 25'd3534751, 25'd1398363, 25'd2485979, 25'd1398363, 25'd3379377, 25'd1631424}}, '{'{-25'd2874413, -25'd971085, 25'd310747, 25'd3806655, -25'd4389306, 25'd2252918, -25'd4622367, 25'd2641352, 25'd1747954}, '{25'd2835570, -25'd4428150, 25'd1670267, 25'd1903328, 25'd2641352, 25'd155374, 25'd3573594, -25'd2641352, 25'd388434}, '{25'd1553737, -25'd3767812, -25'd1709110, -25'd466121, -25'd3806655, 25'd2058701, 25'd3884342, -25'd3573594, 25'd4933114}, '{-25'd3301691, -25'd699182, 25'd2990943, -25'd3340534, -25'd815712, 25'd2136388, -25'd1514893, 25'd3923185, 25'd2835570}, '{25'd1359520, 25'd1825641, -25'd1825641, 25'd4855427, -25'd4195089, -25'd1126459, 25'd2058701, -25'd1126459, -25'd4311619}, '{-25'd4544680, 25'd504964, -25'd1514893, 25'd4156246, 25'd4855427, 25'd3068630, 25'd893399, 25'd2719039, 25'd194217}, '{25'd2641352, 25'd2252918, 25'd3262847, 25'd4311619, 25'd1514893, -25'd1204146, 25'd4933114, 25'd1087616, -25'd3224004}, '{-25'd3767812, -25'd1320676, -25'd4389306, 25'd1476050, 25'd1786797, 25'd2990943, 25'd738025, 25'd4311619, -25'd738025}, '{25'd854555, 25'd2097545, 25'd2641352, -25'd4505837, 25'd504964, 25'd3767812, 25'd2136388, 25'd233061, 25'd155374}}},
    '{'{'{-25'd849103, -25'd3598579, 25'd3355978, -25'd970403, -25'd1051270, 25'd3355978, 25'd4083781, -25'd2345142, -25'd242601}, '{-25'd4488116, -25'd3679446, 25'd3194244, -25'd2830343, -25'd606502, 25'd1051270, 25'd3558146, 25'd2628176, 25'd970403}, '{-25'd2911210, -25'd4649850, 25'd2142974, -25'd1253438, -25'd2709043, 25'd3355978, -25'd3477279, -25'd40433, 25'd4568983}, '{25'd2223841, 25'd4124214, 25'd3275111, -25'd404335, 25'd2628176, 25'd4245515, 25'd646936, -25'd3194244, 25'd1859940}, '{-25'd4205081, -25'd525635, 25'd3922047, -25'd363901, -25'd2142974, 25'd2021674, -25'd283034, -25'd889536, -25'd3598579}, '{-25'd121300, -25'd2385575, -25'd3355978, -25'd525635, 25'd4892450, 25'd1576905, -25'd687369, 25'd970403, 25'd3517712}, '{-25'd80867, 25'd1455605, 25'd3396412, 25'd1617339, 25'd525635, 25'd3800747, 25'd3679446, 25'd4771150, 25'd4892450}, '{-25'd242601, 25'd2183408, -25'd1253438, 25'd1293871, 25'd5135051, 25'd4568983, 25'd4932884, -25'd2911210, -25'd1496039}, '{-25'd3436845, -25'd404335, -25'd2668609, 25'd2628176, 25'd2142974, -25'd808669, -25'd1576905, -25'd3598579, 25'd1415172}}, '{'{25'd2506875, 25'd2870777, -25'd2992077, 25'd444768, -25'd2951644, -25'd2021674, 25'd4568983, 25'd4852017, -25'd3962480}, '{25'd0, 25'd2789910, -25'd2102541, 25'd929970, -25'd3760313, 25'd444768, 25'd1496039, 25'd4447682, 25'd1940807}, '{25'd2668609, 25'd1455605, -25'd4771150, 25'd3639013, -25'd1415172, -25'd404335, 25'd4083781, 25'd5054184, -25'd1091704}, '{25'd3113378, -25'd2870777, 25'd4568983, -25'd2142974, -25'd3922047, -25'd3639013, -25'd4205081, 25'd849103, -25'd4164648}, '{25'd4164648, 25'd2223841, 25'd4043347, 25'd3032511, 25'd2668609, 25'd1213004, 25'd646936, 25'd2385575, -25'd4366815}, '{-25'd3962480, -25'd2021674, -25'd323468, 25'd2749476, -25'd121300, -25'd3558146, -25'd4690283, 25'd2628176, -25'd2830343}, '{25'd5013751, 25'd4285948, -25'd40433, 25'd0, -25'd3436845, -25'd363901, 25'd3072944, -25'd1900373, -25'd1738639}, '{25'd4245515, -25'd323468, -25'd1536472, 25'd2830343, -25'd1657772, 25'd1617339, -25'd2062107, 25'd4892450, -25'd687369}, '{-25'd4407249, -25'd4528549, -25'd2992077, 25'd3355978, -25'd2466442, -25'd4285948, 25'd5013751, 25'd4649850, -25'd4285948}}, '{'{25'd323468, 25'd4083781, -25'd2062107, 25'd1213004, -25'd3436845, 25'd4285948, 25'd3032511, 25'd4245515, -25'd1940807}, '{25'd4771150, -25'd404335, -25'd4366815, -25'd2102541, 25'd3315545, 25'd2709043, 25'd3072944, -25'd363901, -25'd1172571}, '{-25'd363901, -25'd4326382, -25'd3800747, 25'd3032511, -25'd2385575, -25'd4811583, -25'd1859940, -25'd2506875, -25'd2102541}, '{25'd4609416, -25'd2628176, 25'd1617339, 25'd1334305, 25'd3800747, 25'd2911210, -25'd687369, -25'd1415172, 25'd1738639}, '{-25'd3436845, 25'd4852017, 25'd3962480, 25'd3841180, 25'd3477279, 25'd2385575, -25'd80867, -25'd3153811, -25'd4366815}, '{25'd1334305, -25'd3598579, -25'd2547309, -25'd485202, -25'd3315545, 25'd1415172, 25'd404335, 25'd525635, -25'd4002914}, '{-25'd3558146, 25'd2587742, 25'd1859940, 25'd2749476, 25'd4730716, -25'd3679446, 25'd0, -25'd3153811, -25'd2668609}, '{25'd1091704, 25'd3679446, 25'd363901, 25'd2911210, 25'd3922047, 25'd3922047, 25'd2911210, 25'd4124214, 25'd485202}, '{-25'd727803, -25'd2789910, 25'd2021674, -25'd3436845, 25'd3275111, -25'd80867, 25'd1859940, 25'd3275111, 25'd0}}},
    '{'{'{25'd4210595, -25'd620509, -25'd1595594, 25'd753475, -25'd3767374, -25'd975085, -25'd2526357, 25'd0, -25'd3501442}, '{-25'd5052714, 25'd2526357, -25'd5628901, 25'd2792289, -25'd5673223, -25'd2038814, 25'd1462628, 25'd265932, -25'd5584579}, '{-25'd2570679, 25'd177288, 25'd1152373, -25'd3501442, -25'd2437713, 25'd797797, -25'd2615001, -25'd2747967, 25'd4520849}, '{-25'd1994492, -25'd5673223, -25'd310254, -25'd443221, 25'd4299239, 25'd2437713, 25'd4698137, -25'd3501442, 25'd3368476}, '{25'd1063729, -25'd3235510, 25'd4964070, 25'd5097036, -25'd398898, -25'd1063729, 25'd3944663, 25'd3279832, -25'd2216103}, '{-25'd4121951, -25'd1462628, 25'd4210595, -25'd3279832, -25'd4698137, -25'd2747967, -25'd3856018, -25'd2880933, -25'd1196695}, '{-25'd2570679, -25'd2260425, 25'd3501442, 25'd4033307, 25'd1684238, -25'd4520849, -25'd3013900, -25'd1108051, -25'd310254}, '{-25'd177288, -25'd930763, 25'd1418306, 25'd5141358, -25'd1108051, 25'd1285339, 25'd132966, 25'd4432205, 25'd3944663}, '{25'd310254, -25'd975085, 25'd2482035, -25'd531865, 25'd3146866, -25'd2659323, 25'd3102544, 25'd1684238, -25'd2836611}}, '{'{-25'd2038814, -25'd1595594, -25'd4831104, -25'd3678730, -25'd1196695, -25'd4786782, -25'd1462628, -25'd753475, 25'd2083136}, '{25'd132966, -25'd842119, -25'd3324154, 25'd2925255, -25'd5673223, -25'd4254917, 25'd1506950, -25'd487543, -25'd975085}, '{-25'd3058222, -25'd5584579, -25'd664831, -25'd2482035, 25'd1905848, -25'd1994492, 25'd2526357, -25'd1196695, 25'd3634408}, '{-25'd2615001, -25'd1950170, 25'd1684238, 25'd5185680, -25'd1861526, -25'd1905848, 25'd2615001, -25'd3590086, -25'd2747967}, '{25'd3102544, -25'd3811696, -25'd2304747, 25'd3501442, -25'd3900341, -25'd1241017, 25'd3856018, 25'd3102544, -25'd1595594}, '{-25'd5362968, -25'd5673223, -25'd1418306, 25'd3944663, 25'd797797, -25'd4831104, -25'd3102544, 25'd3368476, -25'd1684238}, '{-25'd3013900, 25'd1108051, -25'd2747967, 25'd2792289, 25'd3678730, 25'd1418306, 25'd4033307, 25'd1373984, 25'd3767374}, '{-25'd4742460, -25'd5673223, 25'd265932, -25'd2083136, -25'd443221, 25'd620509, 25'd2792289, 25'd3146866, -25'd2969577}, '{25'd1861526, -25'd2792289, 25'd4033307, -25'd2526357, -25'd3988985, 25'd1196695, -25'd2171781, 25'd930763, 25'd2393391}}, '{'{25'd4520849, -25'd1196695, -25'd5008392, 25'd3324154, -25'd5141358, 25'd1817204, -25'd797797, -25'd3944663, 25'd3501442}, '{25'd1329662, -25'd4742460, -25'd2526357, -25'd2792289, -25'd5451612, 25'd177288, 25'd1506950, -25'd1063729, -25'd3102544}, '{-25'd1063729, -25'd4166273, -25'd4476527, 25'd2083136, 25'd1418306, 25'd2393391, 25'd2349069, 25'd709153, -25'd2526357}, '{25'd177288, -25'd5673223, -25'd4210595, -25'd1373984, 25'd3856018, -25'd398898, 25'd398898, -25'd1506950, 25'd3324154}, '{-25'd2925255, -25'd3634408, -25'd1994492, -25'd1373984, -25'd1772882, -25'd753475, -25'd4121951, 25'd2127458, 25'd1506950}, '{25'd1551272, -25'd4609493, -25'd2615001, -25'd1196695, 25'd1152373, 25'd1728560, 25'd4432205, 25'd1595594, 25'd3900341}, '{-25'd2437713, -25'd398898, 25'd3988985, 25'd975085, -25'd664831, 25'd753475, 25'd310254, 25'd1817204, -25'd265932}, '{-25'd3900341, -25'd5673223, 25'd3102544, 25'd2969577, 25'd1373984, 25'd2304747, -25'd3811696, -25'd4432205, 25'd1905848}, '{-25'd1418306, 25'd177288, 25'd797797, -25'd797797, -25'd2437713, 25'd2083136, 25'd4698137, -25'd3545764, 25'd3634408}}},
    '{'{'{-25'd4136688, -25'd1750137, -25'd318207, -25'd3182068, 25'd1431931, 25'd238655, -25'd3380947, 25'd278431, -25'd2784309}, '{25'd676189, 25'd2346775, -25'd2545654, 25'd2306999, -25'd3341171, -25'd4335567, -25'd4335567, 25'd3818481, 25'd835293}, '{-25'd1153500, 25'd198879, -25'd2585430, -25'd3540051, 25'd4375343, 25'd1073948, -25'd3142292, 25'd2227448, -25'd278431}, '{-25'd556862, 25'd3977585, -25'd3062740, 25'd4256016, 25'd4375343, 25'd3142292, 25'd4057137, -25'd4057137, -25'd3420723}, '{-25'd4653774, 25'd4733326, -25'd1034172, 25'd4892429, -25'd397758, 25'd357983, 25'd3102516, -25'd2426327, 25'd1909241}, '{25'd715965, 25'd3420723, 25'd3341171, -25'd1949017, 25'd914845, 25'd4852654, -25'd1312603, 25'd198879, 25'd4057137}, '{-25'd2028568, -25'd1789913, 25'd3022964, -25'd4057137, 25'd437534, -25'd1591034, -25'd3738930, 25'd437534, 25'd4773102}, '{25'd39776, 25'd4534447, 25'd4892429, 25'd1750137, 25'd1670586, -25'd2108120, -25'd3699154, -25'd954620, 25'd1471706}, '{-25'd517086, 25'd1073948, -25'd1431931, -25'd2863861, 25'd4613998, -25'd4096912, -25'd3738930, -25'd3261620, 25'd1949017}}, '{'{-25'd2346775, 25'd79552, -25'd4653774, -25'd2863861, 25'd4256016, 25'd3380947, -25'd2426327, -25'd3540051, -25'd2426327}, '{25'd3818481, -25'd954620, 25'd596638, 25'd2943413, -25'd4494671, -25'd1591034, -25'd4574223, 25'd119328, 25'd2585430}, '{-25'd3858257, -25'd1670586, -25'd1312603, -25'd119328, -25'd3380947, 25'd3301395, -25'd2824085, -25'd477310, -25'd3977585}, '{25'd1352379, 25'd3858257, 25'd477310, -25'd3182068, -25'd2108120, 25'd2983189, 25'd1551258, 25'd3898033, -25'd1630810}, '{-25'd1312603, 25'd3977585, 25'd278431, 25'd1352379, -25'd1591034, 25'd1630810, -25'd2983189, -25'd2943413, 25'd2625206}, '{25'd0, 25'd1829689, -25'd1153500, 25'd3579826, -25'd1630810, 25'd3858257, 25'd676189, 25'd1789913, -25'd1153500}, '{-25'd1113724, -25'd3858257, -25'd3182068, -25'd636414, -25'd2505878, -25'd715965, 25'd3738930, -25'd119328, -25'd4773102}, '{25'd2545654, -25'd278431, -25'd1750137, 25'd1073948, 25'd278431, -25'd2227448, 25'd159103, 25'd2943413, -25'd3221844}, '{-25'd1392155, 25'd3579826, 25'd4574223, -25'd4256016, 25'd3540051, 25'd1113724, 25'd1591034, -25'd1233051, -25'd3102516}}, '{'{-25'd914845, 25'd3102516, -25'd4494671, -25'd4057137, 25'd1630810, 25'd3500275, 25'd437534, -25'd2664982, 25'd2744534}, '{25'd1471706, -25'd2187672, 25'd119328, -25'd875069, 25'd3380947, -25'd4057137, 25'd914845, 25'd2028568, 25'd3102516}, '{-25'd3142292, 25'd1034172, 25'd3579826, 25'd2068344, 25'd5051533, 25'd2983189, 25'd2426327, -25'd4494671, 25'd1630810}, '{-25'd676189, -25'd715965, 25'd1511482, 25'd4971981, 25'd1949017, -25'd2784309, 25'd1471706, 25'd914845, 25'd3102516}, '{-25'd357983, -25'd2386551, 25'd2585430, 25'd1034172, -25'd477310, 25'd4892429, -25'd1909241, -25'd2306999, 25'd4295792}, '{25'd3420723, 25'd2187672, -25'd2903637, 25'd278431, 25'd278431, -25'd4415119, -25'd3738930, 25'd2943413, 25'd1829689}, '{-25'd1193275, 25'd4057137, -25'd3778706, -25'd1988792, 25'd954620, 25'd4574223, 25'd795517, -25'd994396, 25'd318207}, '{25'd477310, 25'd278431, 25'd2585430, -25'd4335567, -25'd1750137, 25'd4375343, -25'd3540051, 25'd2983189, -25'd3182068}, '{-25'd2784309, -25'd914845, 25'd198879, 25'd3619602, 25'd278431, -25'd2505878, -25'd3699154, -25'd3898033, -25'd2386551}}},
    '{'{'{-25'd2442770, 25'd904729, -25'd4161756, 25'd4433174, -25'd2533242, -25'd4795066, -25'd995202, -25'd3437972, -25'd6514052}, '{-25'd1990405, -25'd3166553, 25'd2352297, -25'd542838, -25'd995202, -25'd5971214, -25'd6152160, -25'd995202, -25'd5156958}, '{-25'd2985607, 25'd3890337, -25'd633311, 25'd5609323, 25'd6604525, -25'd6061687, -25'd3618918, -25'd7509255, -25'd1266621}, '{25'd1628513, -25'd2623715, 25'd1718986, 25'd7328309, 25'd8233038, -25'd11218645, -25'd6152160, -25'd2261824, -25'd4523647}, '{25'd452365, -25'd452365, 25'd5337904, 25'd1447567, 25'd1266621, -25'd7599727, -25'd6604525, 25'd542838, -25'd723784}, '{-25'd3618918, -25'd4704593, 25'd1990405, -25'd2533242, 25'd271419, -25'd5518850, 25'd271419, 25'd1538040, 25'd1085675}, '{-25'd4433174, 25'd1085675, 25'd5247431, 25'd2442770, -25'd90473, -25'd4071283, -25'd7056890, -25'd2080878, -25'd1809459}, '{25'd1718986, 25'd3437972, 25'd4071283, -25'd3076080, 25'd2171351, -25'd9047295, -25'd1899932, -25'd1718986, -25'd4885539}, '{25'd2080878, 25'd2804661, -25'd3166553, -25'd3257026, 25'd0, -25'd8775876, -25'd3347499, -25'd7418782, -25'd1176148}}, '{'{25'd1538040, -25'd1357094, 25'd4523647, 25'd6333106, 25'd1809459, -25'd5880741, -25'd1266621, -25'd6785471, -25'd4252228}, '{25'd3257026, -25'd2985607, 25'd5247431, 25'd2080878, 25'd2261824, -25'd8142565, -25'd7237836, -25'd542838, -25'd7328309}, '{-25'd542838, 25'd4071283, 25'd5247431, 25'd3437972, 25'd4252228, -25'd11580537, -25'd2352297, -25'd6152160, -25'd4795066}, '{-25'd1357094, -25'd995202, 25'd452365, -25'd271419, 25'd6785471, -25'd5156958, -25'd4433174, -25'd5337904, -25'd6966417}, '{25'd3437972, 25'd1447567, 25'd2895134, -25'd180946, 25'd6423579, -25'd6785471, -25'd1266621, -25'd2623715, -25'd452365}, '{25'd904729, -25'd1899932, 25'd4071283, -25'd271419, 25'd2171351, -25'd4523647, -25'd3347499, -25'd2895134, -25'd1809459}, '{-25'd2442770, 25'd361892, -25'd1899932, 25'd1085675, 25'd5428377, -25'd4795066, -25'd271419, -25'd2171351, 25'd180946}, '{-25'd2533242, 25'd1718986, 25'd2261824, 25'd3166553, 25'd1718986, -25'd2352297, -25'd723784, 25'd271419, -25'd361892}, '{25'd3980810, 25'd2533242, 25'd542838, 25'd0, 25'd4523647, -25'd7509255, 25'd1357094, 25'd1357094, -25'd5790269}}, '{'{-25'd3437972, -25'd2171351, 25'd633311, -25'd2261824, 25'd3799864, -25'd10856754, -25'd4704593, -25'd4795066, -25'd4433174}, '{-25'd904729, -25'd361892, 25'd3257026, -25'd1718986, 25'd6152160, -25'd7961619, -25'd7237836, -25'd3166553, -25'd5880741}, '{-25'd4704593, 25'd3257026, 25'd1085675, 25'd6061687, 25'd814257, -25'd8866349, -25'd452365, -25'd1990405, -25'd7599727}, '{25'd1176148, -25'd2352297, 25'd2985607, 25'd5428377, 25'd6694998, -25'd8142565, -25'd4976012, -25'd723784, -25'd5971214}, '{-25'd2352297, 25'd5971214, 25'd1447567, 25'd814257, 25'd271419, -25'd10856754, -25'd2714188, 25'd271419, -25'd6423579}, '{25'd2261824, -25'd3166553, 25'd3166553, 25'd2895134, -25'd814257, -25'd7871146, -25'd7147363, -25'd1266621, -25'd542838}, '{25'd2895134, -25'd1266621, 25'd2714188, -25'd1357094, 25'd180946, -25'd10223443, -25'd7147363, 25'd1447567, -25'd814257}, '{25'd361892, -25'd3257026, -25'd542838, 25'd5699796, 25'd7056890, -25'd6875944, -25'd5066485, -25'd4252228, -25'd3257026}, '{-25'd2804661, -25'd2804661, 25'd5428377, 25'd4704593, 25'd5428377, -25'd4885539, 25'd1176148, -25'd4614120, 25'd361892}}},
    '{'{'{25'd4972365, 25'd844364, 25'd4878546, -25'd4597092, 25'd2486182, -25'd328364, 25'd3377455, 25'd3002182, 25'd4456364}, '{25'd4128001, -25'd2486182, 25'd797455, -25'd234545, -25'd1970182, -25'd2157819, 25'd3799637, 25'd4362546, 25'd4128001}, '{25'd2251637, -25'd3518182, -25'd4362546, -25'd2439273, -25'd1735637, -25'd1641818, 25'd4503274, 25'd328364, 25'd1735637}, '{25'd3612001, -25'd328364, -25'd1688728, 25'd469091, 25'd2204728, -25'd2251637, 25'd1313455, 25'd2626910, -25'd2439273}, '{25'd4644001, -25'd3096001, 25'd1313455, -25'd3189819, 25'd5535274, 25'd1923273, 25'd5863637, 25'd3893455, 25'd985091}, '{-25'd4690910, -25'd281455, -25'd703636, -25'd3846546, -25'd140727, 25'd891273, -25'd4221819, 25'd2110909, 25'd4268728}, '{25'd187636, -25'd4878546, 25'd1172727, -25'd3612001, -25'd4221819, -25'd5347637, -25'd2908364, -25'd1032000, -25'd4081092}, '{-25'd4878546, 25'd891273, -25'd703636, -25'd140727, -25'd1782546, -25'd3189819, 25'd281455, 25'd1078909, 25'd3471273}, '{25'd187636, -25'd4690910, -25'd1970182, 25'd3283637, -25'd3612001, 25'd938182, 25'd0, -25'd3752728, -25'd891273}}, '{'{-25'd2767637, -25'd3846546, -25'd3752728, 25'd3940364, -25'd328364, 25'd891273, -25'd2392364, 25'd844364, -25'd938182}, '{25'd703636, -25'd2345455, -25'd3142910, 25'd2110909, -25'd2110909, -25'd2580000, 25'd1454182, -25'd1548000, 25'd3096001}, '{25'd4221819, -25'd2345455, 25'd4362546, 25'd562909, -25'd4034183, 25'd4644001, -25'd2251637, 25'd2955273, -25'd140727}, '{25'd4456364, -25'd3377455, -25'd1454182, 25'd2580000, 25'd3893455, -25'd281455, -25'd1548000, 25'd2908364, -25'd1360364}, '{25'd4174910, 25'd4409455, -25'd1407273, -25'd2064000, -25'd562909, 25'd703636, -25'd3236728, -25'd3705819, 25'd4690910}, '{-25'd422182, 25'd562909, -25'd4644001, -25'd1782546, -25'd3283637, 25'd3658910, 25'd1032000, -25'd3236728, 25'd4784728}, '{-25'd6004365, -25'd2345455, 25'd46909, -25'd5347637, -25'd1313455, -25'd1219637, -25'd2486182, -25'd5347637, 25'd2908364}, '{25'd1125818, -25'd4784728, -25'd5066183, -25'd140727, -25'd891273, -25'd1313455, 25'd4878546, 25'd1125818, -25'd1829455}, '{-25'd5019274, -25'd4690910, -25'd3002182, -25'd3236728, -25'd93818, 25'd1641818, 25'd4268728, 25'd2298546, 25'd4034183}}, '{'{25'd1313455, 25'd1360364, 25'd234545, 25'd4081092, -25'd46909, 25'd656727, -25'd1923273, 25'd5206910, -25'd187636}, '{25'd3518182, -25'd3893455, -25'd938182, 25'd1548000, -25'd3330546, 25'd1454182, -25'd2861455, 25'd93818, 25'd5253819}, '{25'd4878546, -25'd3799637, -25'd1501091, 25'd2064000, -25'd3330546, -25'd4081092, -25'd3471273, 25'd2345455, 25'd4878546}, '{25'd4972365, -25'd1688728, 25'd4268728, 25'd1501091, 25'd422182, -25'd3236728, 25'd234545, -25'd562909, 25'd1923273}, '{-25'd844364, -25'd4034183, -25'd3940364, 25'd1313455, -25'd656727, -25'd1360364, 25'd4081092, 25'd562909, -25'd1032000}, '{25'd3846546, -25'd234545, 25'd4034183, 25'd3987273, -25'd4034183, 25'd2392364, 25'd938182, -25'd4737819, -25'd2814546}, '{-25'd2580000, 25'd187636, 25'd2204728, -25'd5253819, 25'd375273, 25'd2814546, -25'd4784728, -25'd2673819, 25'd750546}, '{25'd3799637, -25'd3283637, 25'd1032000, 25'd375273, 25'd2345455, 25'd2767637, -25'd2110909, -25'd4081092, -25'd4503274}, '{-25'd3940364, 25'd1594909, -25'd5863637, -25'd5910547, 25'd2767637, 25'd3752728, -25'd3424364, -25'd469091, -25'd1172727}}},
    '{'{'{-25'd2006214, 25'd793154, 25'd3079305, 25'd3219273, 25'd4618957, 25'd1073091, 25'd606530, 25'd1446340, 25'd4385677}, '{25'd2192838, -25'd4572301, -25'd1492996, 25'd3219273, -25'd5038862, -25'd186625, 25'd3965771, -25'd4105740, 25'd4572301}, '{-25'd3079305, 25'd4432333, 25'd2706056, -25'd2939336, -25'd559874, -25'd2332807, -25'd2846024, -25'd4525645, 25'd2566087}, '{-25'd3265929, -25'd3825803, -25'd2985993, -25'd2519431, 25'd2332807, 25'd2939336, 25'd839810, 25'd4665613, 25'd4152396}, '{25'd793154, 25'd1679621, 25'd2612743, -25'd2006214, -25'd5785361, -25'd1492996, 25'd746498, 25'd3125961, -25'd4245708}, '{25'd2659400, 25'd3452554, 25'd979779, -25'd5645392, -25'd4292364, 25'd139968, 25'd979779, -25'd1632965, 25'd1726277}, '{25'd1819589, -25'd2846024, -25'd1726277, 25'd2472775, -25'd4199052, -25'd4898894, -25'd3219273, 25'd2379463, 25'd979779}, '{25'd4339020, -25'd3639178, 25'd2052870, 25'd793154, 25'd186625, -25'd1446340, 25'd1353028, -25'd4618957, 25'd2706056}, '{-25'd3219273, -25'd2892680, 25'd5038862, 25'd746498, 25'd1306372, -25'd2846024, 25'd4292364, 25'd2892680, -25'd5085519}}, '{'{-25'd186625, -25'd2426119, -25'd1166403, 25'd4852238, 25'd1306372, -25'd1866245, -25'd2239494, 25'd3219273, -25'd2892680}, '{-25'd4618957, 25'd2472775, 25'd933123, -25'd1306372, -25'd3685835, 25'd1306372, -25'd653186, 25'd326593, 25'd793154}, '{25'd4385677, 25'd2892680, 25'd2146182, 25'd3032649, 25'd1632965, -25'd2146182, 25'd3405898, 25'd3452554, 25'd3079305}, '{-25'd3405898, -25'd373249, 25'd1866245, -25'd4525645, 25'd933123, 25'd793154, -25'd1259716, 25'd2846024, -25'd1866245}, '{25'd5132175, -25'd3732491, -25'd2892680, 25'd3452554, -25'd3779147, -25'd839810, -25'd1213059, -25'd1213059, 25'd5318799}, '{25'd2286151, -25'd3405898, 25'd1213059, -25'd2985993, -25'd5971985, -25'd5365455, 25'd746498, 25'd4618957, -25'd1632965}, '{25'd4432333, 25'd3825803, 25'd2052870, -25'd1539652, -25'd2426119, -25'd886467, -25'd2612743, 25'd4012427, -25'd2985993}, '{25'd4478989, 25'd93312, -25'd886467, -25'd4292364, -25'd3079305, -25'd3032649, 25'd3592522, 25'd4245708, -25'd933123}, '{-25'd559874, 25'd1819589, -25'd3639178, 25'd4618957, 25'd886467, -25'd1399684, 25'd606530, 25'd2519431, -25'd2659400}}, '{'{-25'd3312585, 25'd2006214, -25'd2239494, 25'd1632965, -25'd93312, 25'd1026435, -25'd1353028, 25'd1772933, 25'd559874}, '{-25'd2566087, 25'd3779147, -25'd326593, -25'd2706056, -25'd1679621, -25'd653186, -25'd1819589, 25'd2472775, -25'd2939336}, '{25'd3359242, 25'd839810, 25'd1259716, 25'd373249, 25'd3872459, -25'd5178831, -25'd3732491, -25'd1819589, 25'd4292364}, '{-25'd2752712, 25'd2286151, 25'd1772933, -25'd3545866, -25'd5598736, 25'd139968, -25'd4618957, 25'd4245708, -25'd839810}, '{-25'd419905, 25'd3265929, -25'd2892680, -25'd3592522, 25'd3359242, -25'd2892680, 25'd886467, -25'd2612743, 25'd4385677}, '{25'd2659400, 25'd2146182, -25'd4245708, -25'd3965771, -25'd3452554, -25'd4199052, 25'd886467, 25'd2706056, 25'd5365455}, '{25'd1539652, -25'd513217, 25'd1446340, -25'd746498, -25'd5272143, -25'd3172617, -25'd1772933, 25'd4478989, 25'd2286151}, '{25'd4945550, 25'd2286151, 25'd3452554, -25'd3779147, 25'd93312, 25'd1213059, -25'd2286151, -25'd1632965, 25'd2939336}, '{25'd5178831, 25'd46656, -25'd2799368, -25'd2706056, -25'd3499210, 25'd2379463, -25'd1213059, 25'd1866245, -25'd326593}}},
    '{'{'{-25'd2564129, -25'd3025673, 25'd205130, 25'd307696, 25'd923087, 25'd3692346, -25'd2410282, -25'd2923107, -25'd3538498}, '{-25'd3025673, -25'd2871825, -25'd4820563, 25'd153848, -25'd4717998, 25'd2974390, -25'd1025652, -25'd2564129, -25'd4307737}, '{-25'd3487216, -25'd3641064, 25'd1743608, 25'd1538478, 25'd1230782, 25'd1487195, 25'd3435933, 25'd3282086, -25'd5487237}, '{-25'd2153869, 25'd1589760, -25'd974369, -25'd2102586, 25'd3230803, -25'd2512847, 25'd1487195, 25'd4871846, -25'd871804}, '{-25'd769239, -25'd3333368, -25'd3282086, 25'd6102628, -25'd2410282, 25'd2666694, -25'd1948738, 25'd1794891, 25'd461543}, '{-25'd1692325, 25'd564108, 25'd102565, 25'd1538478, 25'd2871825, -25'd1282065, -25'd358978, -25'd1076934, 25'd1846173}, '{-25'd4153889, -25'd3846194, 25'd410261, 25'd153848, 25'd1897456, -25'd3794911, 25'd769239, -25'd615391, -25'd3230803}, '{25'd4307737, 25'd4153889, 25'd4717998, 25'd4000042, -25'd871804, -25'd1641043, 25'd4615433, 25'd3538498, 25'd2615412}, '{-25'd1487195, -25'd1641043, -25'd1692325, -25'd2512847, -25'd4359020, 25'd1897456, -25'd3538498, -25'd2461564, -25'd2820542}}, '{'{-25'd1076934, -25'd5435954, 25'd3435933, -25'd2051303, 25'd4769281, -25'd3179520, -25'd615391, -25'd512826, 25'd1948738}, '{-25'd2820542, -25'd1641043, 25'd2461564, -25'd615391, -25'd1692325, 25'd307696, 25'd3538498, -25'd5282106, -25'd1794891}, '{25'd871804, -25'd2615412, 25'd2307716, 25'd205130, 25'd1230782, 25'd4820563, 25'd2256434, -25'd1179499, -25'd5282106}, '{-25'd2564129, 25'd2871825, 25'd4769281, 25'd1589760, -25'd923087, 25'd4102607, 25'd1179499, 25'd2512847, -25'd2974390}, '{25'd2461564, -25'd1487195, 25'd6512888, 25'd1487195, 25'd3897477, 25'd3794911, 25'd1846173, -25'd3948759, -25'd2307716}, '{25'd3282086, -25'd1435912, 25'd974369, -25'd1743608, -25'd2358999, 25'd153848, 25'd0, -25'd4307737, 25'd1948738}, '{-25'd923087, -25'd3076955, -25'd564108, -25'd358978, 25'd5641084, 25'd5179541, 25'd3641064, -25'd2564129, 25'd1846173}, '{-25'd1897456, -25'd410261, 25'd5641084, -25'd3025673, 25'd4717998, 25'd4666715, 25'd3589781, 25'd1179499, 25'd2717977}, '{-25'd256413, -25'd205130, 25'd615391, 25'd2512847, 25'd3641064, -25'd3948759, 25'd1794891, 25'd3128238, -25'd2000021}}, '{'{25'd3076955, 25'd410261, -25'd4512868, 25'd4923128, -25'd2615412, -25'd2461564, -25'd3025673, 25'd3743629, -25'd5487237}, '{25'd2358999, 25'd2871825, 25'd3743629, -25'd1641043, 25'd1128217, 25'd871804, -25'd3897477, -25'd769239, 25'd1435912}, '{-25'd4410302, -25'd4974411, 25'd2769260, 25'd769239, 25'd1230782, 25'd2923107, 25'd0, -25'd4820563, -25'd102565}, '{25'd2000021, -25'd3589781, 25'd1743608, -25'd1179499, 25'd5743650, 25'd1641043, -25'd2205151, 25'd1025652, 25'd3333368}, '{-25'd923087, -25'd2461564, 25'd1692325, 25'd2820542, -25'd1487195, 25'd3282086, 25'd2717977, 25'd3487216, -25'd1128217}, '{-25'd871804, -25'd4359020, -25'd512826, 25'd4820563, 25'd1025652, 25'd2871825, 25'd5846215, 25'd5230824, 25'd1846173}, '{-25'd3076955, -25'd1025652, 25'd2102586, 25'd1589760, 25'd3025673, 25'd923087, -25'd871804, 25'd1487195, 25'd3641064}, '{25'd2666694, -25'd307696, 25'd923087, 25'd4666715, -25'd2820542, -25'd1641043, 25'd4153889, -25'd3948759, 25'd2256434}, '{25'd153848, -25'd3179520, -25'd4153889, 25'd1025652, -25'd2974390, 25'd2410282, 25'd3538498, 25'd2153869, -25'd4769281}}},
    '{'{'{-25'd4132229, -25'd1186917, 25'd4308068, -25'd351679, 25'd219799, -25'd1582556, 25'd219799, -25'd3736590, 25'd1055037}, '{-25'd5275186, -25'd527519, -25'd2505713, -25'd2989272, -25'd1758395, -25'd1846315, 25'd351679, 25'd3648670, 25'd3956389}, '{-25'd615438, 25'd1055037, 25'd4044309, -25'd1538596, -25'd5538945, -25'd923157, 25'd1406716, 25'd1406716, 25'd2637593}, '{25'd3824510, 25'd2505713, 25'd1318796, 25'd703358, -25'd2461753, -25'd2945312, -25'd4483908, -25'd4439948, -25'd483559}, '{25'd4088269, 25'd3121151, 25'd3648670, -25'd1406716, -25'd263759, 25'd175840, -25'd4044309, 25'd3824510, 25'd3253031}, '{-25'd3868469, -25'd2901352, -25'd5363105, -25'd5626865, 25'd1670475, -25'd1978195, -25'd615438, 25'd659398, -25'd1670475}, '{25'd4747667, 25'd3604710, -25'd2461753, -25'd2154034, -25'd4615787, -25'd1758395, 25'd131880, -25'd2373833, 25'd1362756}, '{25'd483559, 25'd1538596, -25'd3165111, 25'd2505713, -25'd527519, -25'd1450676, 25'd483559, -25'd2154034, 25'd1846315}, '{25'd3077192, 25'd4264108, 25'd1318796, -25'd3692630, 25'd3253031, -25'd2725513, 25'd3780550, -25'd4044309, -25'd4791627}}, '{'{25'd2417793, 25'd659398, 25'd483559, -25'd3209071, 25'd747318, 25'd3340951, 25'd4527868, 25'd1230877, 25'd2241954}, '{25'd3165111, 25'd4395988, -25'd2285914, 25'd3868469, 25'd1142957, 25'd4352028, -25'd3296991, -25'd2373833, 25'd4967466}, '{25'd219799, -25'd615438, 25'd3384911, 25'd4308068, 25'd175840, -25'd175840, 25'd87920, 25'd131880, 25'd4967466}, '{25'd351679, -25'd1934235, 25'd3033232, 25'd1230877, 25'd1274837, -25'd2285914, -25'd1802355, 25'd3560750, 25'd4000349}, '{-25'd4308068, -25'd1055037, 25'd3296991, 25'd1230877, -25'd2329874, 25'd1758395, 25'd2461753, 25'd2285914, 25'd2813432}, '{-25'd1978195, 25'd1186917, 25'd2461753, 25'd879198, 25'd2857392, 25'd263759, 25'd2154034, 25'd483559, 25'd1362756}, '{-25'd43960, 25'd1098997, 25'd4571827, -25'd3472830, 25'd3209071, -25'd2241954, 25'd571478, -25'd3296991, -25'd2505713}, '{-25'd3077192, 25'd4000349, 25'd1055037, 25'd483559, -25'd2022154, 25'd3472830, 25'd2637593, -25'd483559, -25'd2725513}, '{25'd2066114, 25'd4395988, 25'd1142957, 25'd2945312, -25'd2241954, -25'd1230877, -25'd1098997, -25'd3516790, 25'd3340951}}, '{'{25'd3253031, 25'd2022154, -25'd1055037, 25'd1318796, 25'd307719, 25'd1450676, -25'd5451025, -25'd571478, -25'd571478}, '{-25'd4308068, 25'd1318796, -25'd4483908, -25'd1406716, -25'd1934235, 25'd2154034, 25'd439599, 25'd1055037, 25'd4088269}, '{25'd4000349, 25'd2373833, 25'd967117, -25'd4967466, -25'd175840, -25'd483559, 25'd1890275, -25'd2813432, -25'd3604710}, '{-25'd4791627, -25'd219799, 25'd3165111, 25'd1802355, 25'd1538596, -25'd835238, -25'd2110074, 25'd2197994, 25'd4747667}, '{25'd4308068, -25'd2066114, -25'd1011077, -25'd1758395, -25'd4571827, -25'd3253031, -25'd3560750, -25'd3736590, -25'd4483908}, '{-25'd527519, 25'd791278, -25'd2066114, -25'd5011426, 25'd1142957, -25'd2593633, 25'd1802355, -25'd1978195, 25'd1714435}, '{25'd2329874, -25'd4527868, 25'd1582556, -25'd3077192, -25'd4395988, -25'd5275186, 25'd4483908, -25'd3868469, 25'd1011077}, '{25'd2241954, 25'd3296991, -25'd4747667, -25'd43960, 25'd1098997, 25'd2329874, -25'd1582556, -25'd1846315, -25'd2461753}, '{-25'd1978195, -25'd5319145, 25'd4439948, -25'd2110074, -25'd1142957, -25'd87920, 25'd1582556, 25'd967117, 25'd3033232}}},
    '{'{'{-25'd1526025, -25'd1017350, -25'd626061, -25'd3404209, 25'd1134736, -25'd978221, 25'd4695461, 25'd1604282, 25'd2699890}, '{-25'd4734589, -25'd1604282, 25'd3365080, -25'd4734589, -25'd626061, -25'd1408638, -25'd2034700, 25'd3756368, -25'd39129}, '{-25'd2778148, -25'd626061, 25'd1878184, -25'd508675, 25'd1095607, -25'd2386859, -25'd3286822, -25'd2112957, -25'd1173865}, '{25'd3325951, -25'd4695461, -25'd430417, 25'd2269473, 25'd1760798, -25'd547804, 25'd4656332, 25'd4734589, 25'd2191215}, '{-25'd3012921, 25'd352160, 25'd2230344, 25'd4147657, -25'd4578074, 25'd3404209, -25'd782577, 25'd3130307, -25'd2934663}, '{25'd3756368, -25'd3756368, 25'd4499816, -25'd3012921, 25'd3247694, 25'd430417, 25'd4069399, 25'd4460688, -25'd2739019}, '{25'd3247694, 25'd3286822, 25'd4225915, 25'd1643411, -25'd469546, 25'd3521595, -25'd234773, 25'd4421559, -25'd1878184}, '{25'd4617203, -25'd2895534, -25'd4538945, -25'd2778148, 25'd3482467, -25'd2073828, -25'd1760798, 25'd978221, -25'd2856405}, '{-25'd4812847, 25'd3169436, 25'd782577, -25'd2973792, -25'd78258, -25'd2152086, -25'd2543374, 25'd1486896, 25'd2269473}}, '{'{25'd2973792, 25'd1995571, -25'd391288, -25'd273902, -25'd3208565, 25'd1056479, 25'd2660761, -25'd4656332, -25'd1604282}, '{25'd665190, -25'd1017350, -25'd782577, 25'd3443338, -25'd430417, 25'd2425988, -25'd4343301, -25'd352160, 25'd1408638}, '{25'd3952013, -25'd3443338, -25'd1095607, -25'd2073828, -25'd5008491, 25'd4773718, -25'd39129, -25'd3991141, -25'd156515}, '{25'd1369509, 25'd3521595, 25'd1134736, -25'd4538945, -25'd4343301, 25'd156515, 25'd2073828, 25'd3247694, 25'd2699890}, '{-25'd2660761, 25'd2621632, 25'd1760798, -25'd4891105, 25'd4069399, 25'd2112957, -25'd1526025, -25'd1917313, 25'd352160}, '{-25'd4812847, 25'd4225915, 25'd1799927, -25'd1995571, 25'd1565154, -25'd1330380, 25'd743448, 25'd352160, 25'd2191215}, '{25'd1134736, 25'd4147657, -25'd3012921, 25'd3834626, -25'd1682540, 25'd2347730, 25'd3091178, 25'd2191215, -25'd1878184}, '{25'd626061, 25'd3404209, -25'd2934663, 25'd2425988, -25'd3482467, 25'd4304172, -25'd860834, -25'd2817276, -25'd3208565}, '{-25'd3169436, -25'd3404209, -25'd1995571, 25'd2504246, 25'd2073828, 25'd3286822, -25'd2269473, -25'd2817276, -25'd1956442}}, '{'{-25'd626061, 25'd3599853, -25'd2112957, -25'd4734589, 25'd4460688, 25'd743448, -25'd2386859, -25'd3638982, -25'd234773}, '{25'd1760798, 25'd4304172, 25'd1565154, 25'd273902, -25'd3834626, 25'd3365080, 25'd4147657, -25'd1956442, 25'd2582503}, '{25'd1447767, 25'd3678111, 25'd1682540, 25'd313031, -25'd156515, -25'd78258, 25'd2425988, 25'd3286822, -25'd2895534}, '{-25'd899963, 25'd1956442, -25'd4225915, 25'd4617203, 25'd4382430, 25'd2465117, -25'd1212994, -25'd3208565, -25'd1095607}, '{-25'd1839055, 25'd939092, 25'd1799927, -25'd156515, -25'd1212994, 25'd3795497, 25'd704319, -25'd1212994, 25'd1095607}, '{25'd782577, -25'd4382430, 25'd3443338, -25'd1799927, -25'd2230344, 25'd1095607, 25'd117387, 25'd3834626, 25'd1369509}, '{-25'd1252123, 25'd4969362, -25'd3169436, 25'd2817276, -25'd273902, 25'd3012921, 25'd3325951, 25'd3599853, -25'd1799927}, '{-25'd117387, -25'd3091178, -25'd391288, -25'd234773, -25'd4382430, 25'd626061, -25'd78258, 25'd1839055, -25'd4186786}, '{-25'd939092, 25'd3247694, -25'd352160, 25'd1721669, 25'd2543374, -25'd2621632, 25'd1095607, 25'd2152086, -25'd939092}}},
    '{'{'{-25'd3438176, 25'd2115801, -25'd2569187, -25'd3362612, 25'd2833662, -25'd2304712, 25'd2758098, -25'd1435722, 25'd2682533}, '{-25'd1473504, -25'd3249266, 25'd453386, 25'd4269384, -25'd604515, 25'd2153583, 25'd755643, 25'd604515, -25'd2304712}, '{25'd1813544, 25'd1360158, -25'd1926890, -25'd264475, 25'd4193820, -25'd680079, -25'd264475, -25'd2229147, 25'd3438176}, '{25'd2115801, -25'd604515, -25'd3702651, 25'd2833662, -25'd3853780, 25'd0, 25'd1020118, -25'd2266929, -25'd2569187}, '{25'd377822, 25'd944554, 25'd1851326, -25'd3324830, 25'd4118255, -25'd566732, 25'd4118255, 25'd2795880, 25'd3211483}, '{-25'd1322376, -25'd491168, -25'd3702651, 25'd1813544, 25'd2380276, -25'd1549068, 25'd1435722, -25'd1360158, -25'd3589305}, '{-25'd2531405, 25'd2002454, -25'd717861, 25'd3627087, 25'd3815998, -25'd1095683, -25'd1813544, -25'd151129, 25'd1095683}, '{-25'd1624633, -25'd3362612, -25'd1322376, -25'd831207, 25'd4798334, -25'd3362612, 25'd2644751, -25'd3740434, 25'd3098137}, '{-25'd3778216, -25'd1851326, 25'd2984790, -25'd2644751, 25'd113346, -25'd2229147, -25'd4193820, -25'd4684988, -25'd2380276}}, '{'{-25'd4193820, -25'd3513741, 25'd4193820, 25'd944554, -25'd4382730, -25'd4609423, 25'd3249266, 25'd1813544, -25'd75564}, '{-25'd4193820, 25'd831207, -25'd4193820, 25'd3551523, -25'd3287048, -25'd4118255, -25'd755643, -25'd2040237, 25'd3249266}, '{-25'd2115801, 25'd2266929, -25'd2644751, 25'd0, -25'd3475959, -25'd3060355, 25'd3098137, 25'd982336, 25'd264475}, '{25'd1775761, 25'd3475959, 25'd3324830, -25'd3400394, -25'd1209029, -25'd604515, -25'd1057900, 25'd2380276, -25'd1889108}, '{25'd1322376, 25'd4004909, -25'd2644751, -25'd1549068, -25'd4382730, 25'd2342494, -25'd4269384, -25'd1322376, -25'd1586851}, '{25'd2984790, 25'd2531405, -25'd491168, -25'd1775761, 25'd3853780, -25'd4231602, 25'd717861, 25'd4684988, 25'd3664869}, '{-25'd4420512, 25'd3702651, -25'd1322376, -25'd4269384, -25'd1775761, -25'd1813544, 25'd1700197, -25'd755643, -25'd377822}, '{25'd1775761, -25'd2682533, -25'd4307166, 25'd2153583, 25'd2115801, 25'd1133465, 25'd4533859, -25'd4118255, -25'd2153583}, '{25'd2115801, 25'd3287048, -25'd4042691, -25'd4798334, -25'd2531405, -25'd3815998, 25'd340039, 25'd226693, 25'd680079}}, '{'{-25'd3551523, 25'd1397940, 25'd868990, -25'd340039, -25'd4836116, -25'd302257, -25'd906772, 25'd3211483, 25'd793425}, '{25'd4609423, -25'd2078019, 25'd188911, 25'd528950, -25'd37782, 25'd4722770, -25'd1737979, -25'd4231602, -25'd4344948}, '{-25'd831207, 25'd2455840, -25'd2531405, 25'd2833662, 25'd2833662, -25'd642297, 25'd2342494, 25'd4647205, 25'd1360158}, '{25'd3060355, 25'd1851326, 25'd4496077, 25'd188911, -25'd944554, 25'd3249266, 25'd1473504, -25'd3249266, 25'd528950}, '{-25'd2002454, -25'd4684988, -25'd4684988, 25'd2304712, 25'd717861, -25'd2833662, -25'd3475959, -25'd2229147, -25'd4231602}, '{25'd2493622, -25'd1095683, -25'd2229147, -25'd1964672, 25'd4080473, -25'd4722770, 25'd2682533, 25'd0, -25'd2871444}, '{-25'd2002454, 25'd302257, -25'd3324830, -25'd3287048, 25'd0, -25'd3551523, -25'd528950, -25'd415604, 25'd3098137}, '{-25'd4760552, 25'd2569187, -25'd4042691, -25'd642297, 25'd1095683, -25'd4118255, -25'd3060355, -25'd4609423, -25'd1020118}, '{25'd1435722, -25'd3287048, 25'd2984790, 25'd604515, -25'd1397940, 25'd3287048, 25'd1473504, 25'd2531405, -25'd3627087}}},
    '{'{'{25'd4541588, 25'd123861, 25'd4211290, -25'd990892, -25'd1734061, 25'd1445051, 25'd4665449, -25'd2353368, -25'd1156040}, '{25'd123861, -25'd165149, 25'd3591983, 25'd1321189, 25'd4913172, -25'd3096537, 25'd3426834, 25'd2229507, 25'd1899209}, '{25'd2724953, -25'd660595, -25'd206436, 25'd3013963, -25'd2601091, -25'd1486338, 25'd4417726, 25'd1445051, -25'd1362476}, '{-25'd3798419, -25'd1692774, 25'd4871885, -25'd1321189, -25'd1486338, 25'd4170003, -25'd2229507, 25'd784456, 25'd1238615}, '{25'd3633270, -25'd4624162, 25'd412872, -25'd2353368, 25'd3220398, 25'd2807527, -25'd2559804, 25'd990892, 25'd4004854}, '{-25'd578020, 25'd619307, -25'd165149, -25'd1940496, -25'd1238615, 25'd3674557, 25'd4170003, 25'd2105645, 25'd4128716}, '{25'd5078321, -25'd2023071, -25'd123861, -25'd2724953, 25'd4748023, -25'd3261686, 25'd247723, 25'd867030, 25'd784456}, '{25'd3261686, -25'd990892, -25'd2518517, -25'd3426834, 25'd2146932, 25'd4170003, 25'd1527625, 25'd2312081, -25'd2023071}, '{-25'd3880993, 25'd4128716, 25'd1775348, 25'd2394655, 25'd2435942, -25'd3963567, 25'd2312081, 25'd4541588, 25'd536733}}, '{'{25'd1775348, -25'd4376439, -25'd3550696, 25'd949605, 25'd1073466, 25'd2229507, 25'd3055250, -25'd2435942, 25'd1073466}, '{25'd2435942, 25'd1568912, 25'd4871885, 25'd4004854, -25'd990892, -25'd2394655, 25'd4211290, -25'd536733, -25'd4624162}, '{-25'd3013963, -25'd3798419, -25'd619307, 25'd3179111, -25'd2807527, -25'd4376439, -25'd4624162, -25'd4128716, 25'd4789310}, '{-25'd2229507, -25'd4128716, 25'd4541588, 25'd4252577, -25'd1734061, -25'd3096537, -25'd4004854, 25'd3880993, 25'd536733}, '{25'd3798419, 25'd2807527, -25'd82574, -25'd1073466, 25'd1651486, -25'd743169, -25'd2477230, -25'd743169, -25'd1073466}, '{-25'd2312081, -25'd2064358, 25'd4789310, -25'd1527625, 25'd1238615, 25'd1403763, 25'd4624162, -25'd4417726, -25'd1114753}, '{25'd3344260, 25'd82574, -25'd4913172, -25'd4417726, -25'd82574, -25'd3220398, -25'd743169, -25'd3220398, 25'd1692774}, '{-25'd1032179, 25'd4087429, 25'd4417726, -25'd2270794, 25'd1527625, 25'd660595, 25'd908318, 25'd330297, -25'd536733}, '{-25'd2188219, 25'd1568912, 25'd3096537, -25'd3426834, 25'd3509409, -25'd4582875, -25'd2724953, 25'd3468121, 25'd743169}}, '{'{-25'd2848814, 25'd1610199, -25'd3261686, -25'd2518517, 25'd2188219, 25'd1527625, -25'd2518517, 25'd1279902, 25'd5243469}, '{25'd1486338, 25'd4995746, -25'd3013963, 25'd2435942, 25'd495446, 25'd3137824, -25'd1734061, 25'd4541588, 25'd1527625}, '{25'd4748023, -25'd289010, -25'd2312081, 25'd701882, 25'd2188219, 25'd4871885, -25'd1032179, 25'd4335152, -25'd3179111}, '{-25'd1568912, 25'd3757132, 25'd867030, 25'd1321189, -25'd2518517, 25'd3509409, 25'd2559804, 25'd2477230, 25'd1651486}, '{-25'd3715844, -25'd1981784, -25'd1238615, 25'd3509409, 25'd3179111, -25'd2972675, -25'd3509409, 25'd4541588, -25'd3757132}, '{-25'd3013963, -25'd82574, 25'd2766240, 25'd2270794, -25'd4582875, -25'd1527625, -25'd3963567, 25'd1073466, 25'd4830598}, '{-25'd2188219, 25'd1816635, -25'd2477230, 25'd1279902, -25'd2559804, 25'd412872, 25'd908318, 25'd1940496, -25'd3798419}, '{-25'd1568912, 25'd2023071, -25'd82574, 25'd4004854, -25'd371584, 25'd4665449, -25'd908318, 25'd1403763, -25'd3302973}, '{-25'd412872, 25'd5078321, 25'd3922280, -25'd165149, 25'd1734061, 25'd3220398, 25'd2146932, -25'd1403763, -25'd495446}}},
    '{'{'{-25'd2945959, 25'd1568627, -25'd1759923, -25'd2372071, 25'd497370, 25'd3558106, -25'd3175514, 25'd459110, -25'd1339072}, '{-25'd1874701, 25'd1759923, -25'd2372071, 25'd2601626, 25'd459110, -25'd2716403, -25'd2716403, -25'd3481588, 25'd1836442}, '{25'd2639885, 25'd4323290, 25'd3787661, 25'd765184, -25'd459110, -25'd765184, -25'd76518, 25'd4782400, -25'd994739}, '{-25'd4705882, -25'd1300813, 25'd4055476, -25'd4591104, -25'd4820660, 25'd3252032, 25'd4285031, -25'd726925, 25'd1262554}, '{-25'd4782400, -25'd1912960, 25'd1415591, -25'd4629364, 25'd3252032, -25'd535629, 25'd994739, -25'd994739, -25'd1262554}, '{25'd4323290, -25'd2563367, 25'd306074, 25'd2333811, 25'd2525107, -25'd994739, 25'd4744141, -25'd3864180, -25'd650406}, '{-25'd4131994, -25'd2869440, -25'd4017216, -25'd2486848, 25'd1377331, -25'd1836442, -25'd4552845, -25'd2142515, -25'd3060736}, '{-25'd1568627, -25'd459110, -25'd3749402, -25'd2869440, -25'd535629, -25'd4246772, -25'd1683405, -25'd3558106, -25'd191296}, '{25'd841702, 25'd1989479, -25'd4017216, 25'd2792922, -25'd3137255, -25'd191296, -25'd1147776, 25'd726925, 25'd4514586}}, '{'{25'd1568627, 25'd3634624, -25'd459110, -25'd114778, -25'd2831181, -25'd3634624, 25'd1453850, -25'd1912960, -25'd4285031}, '{-25'd2716403, 25'd1224295, 25'd382592, 25'd3481588, -25'd76518, -25'd3098995, 25'd3405069, 25'd4782400, -25'd1606887}, '{-25'd650406, -25'd3864180, -25'd2907699, 25'd4438068, 25'd4705882, -25'd459110, 25'd2333811, 25'd1032998, 25'd3864180}, '{-25'd3290291, -25'd2984218, -25'd2180775, -25'd688666, -25'd1989479, -25'd3711143, 25'd3596365, 25'd2104256, -25'd3825920}, '{25'd1415591, -25'd191296, -25'd2372071, 25'd4017216, -25'd879962, -25'd2372071, -25'd1071258, 25'd4552845, -25'd4591104}, '{25'd2065997, 25'd2448589, -25'd1530368, -25'd4820660, -25'd3252032, -25'd688666, 25'd1453850, 25'd1721664, 25'd3978957}, '{25'd2065997, 25'd153037, -25'd2525107, 25'd3749402, -25'd1262554, -25'd4208512, -25'd1530368, 25'd191296, -25'd1377331}, '{-25'd2563367, -25'd3366810, 25'd3711143, 25'd4170253, 25'd2754663, 25'd1645146, 25'd3672884, 25'd1300813, -25'd3098995}, '{-25'd4897178, -25'd4399808, 25'd1568627, -25'd4055476, -25'd3519847, -25'd1759923, -25'd2563367, 25'd2792922, 25'd2716403}}, '{'{25'd153037, -25'd765184, -25'd2333811, -25'd3749402, 25'd4705882, 25'd2869440, 25'd2984218, -25'd2180775, -25'd2448589}, '{25'd1530368, -25'd1262554, 25'd3366810, 25'd1300813, 25'd1645146, 25'd191296, -25'd2869440, 25'd4285031, -25'd1109517}, '{25'd3252032, -25'd1186035, -25'd1186035, -25'd3443328, 25'd1798183, 25'd3443328, -25'd956480, -25'd4093735, -25'd3787661}, '{-25'd2104256, -25'd3864180, -25'd4858919, -25'd1606887, 25'd2372071, -25'd306074, -25'd3634624, 25'd765184, 25'd2907699}, '{-25'd2448589, 25'd229555, 25'd3022477, 25'd1798183, 25'd1032998, -25'd4820660, -25'd3328551, 25'd3443328, -25'd2486848}, '{-25'd344333, -25'd2372071, 25'd1147776, -25'd1492109, -25'd76518, -25'd4170253, -25'd4820660, -25'd3787661, 25'd2831181}, '{25'd2525107, -25'd4399808, -25'd3596365, 25'd2372071, 25'd3328551, 25'd3137255, 25'd612147, 25'd573888, 25'd1836442}, '{-25'd1798183, -25'd612147, -25'd3634624, -25'd918221, -25'd4399808, 25'd4552845, -25'd3825920, 25'd4399808, 25'd4208512}, '{25'd2372071, -25'd38259, -25'd2372071, -25'd1951219, -25'd1224295, 25'd2792922, -25'd2639885, -25'd3405069, 25'd1415591}}},
    '{'{'{25'd3366118, 25'd990035, 25'd2217678, 25'd3643328, 25'd3762132, -25'd2811699, -25'd1663258, -25'd2613692, -25'd673224}, '{-25'd1821664, 25'd1227643, -25'd3366118, 25'd316811, 25'd1504853, 25'd277210, 25'd2574090, -25'd3960139, -25'd1346447}, '{25'd1188042, -25'd2534489, 25'd1623657, -25'd4514558, -25'd356412, -25'd554419, 25'd1782062, 25'd4158146, 25'd4118544}, '{25'd2059272, -25'd1029636, -25'd1227643, 25'd2970104, 25'd1702860, 25'd4078943, -25'd1940468, 25'd2494887, -25'd4672964}, '{-25'd1029636, -25'd2059272, -25'd2415685, 25'd831629, 25'd0, 25'd4474957, -25'd4910572, -25'd1267244, -25'd1346447}, '{-25'd277210, -25'd1465251, 25'd3286915, -25'd1861265, 25'd1861265, -25'd3762132, 25'd1623657, 25'd3524524, 25'd1584056}, '{-25'd1306846, 25'd4752167, 25'd4791768, 25'd3484922, -25'd4752167, 25'd910832, 25'd2613692, -25'd1702860, 25'd594021}, '{-25'd3722530, -25'd1861265, -25'd2296881, 25'd1227643, -25'd4197747, 25'd514818, 25'd2970104, 25'd4474957, -25'd4831369}, '{25'd2376083, 25'd396014, -25'd4276950, -25'd2217678, 25'd3524524, 25'd2178076, 25'd2376083, 25'd4395754, 25'd1782062}}, '{'{-25'd4237349, 25'd2019671, 25'd2257279, -25'd3128510, 25'd594021, 25'd1544454, 25'd2059272, 25'd3286915, 25'd3405719}, '{25'd3405719, -25'd1623657, 25'd2772097, -25'd3722530, -25'd4039342, -25'd316811, 25'd2534489, 25'd2098874, 25'd4158146}, '{25'd2811699, -25'd2930503, 25'd1386049, 25'd2336482, -25'd4712565, -25'd4989775, -25'd118804, 25'd3128510, -25'd1584056}, '{25'd1821664, -25'd237608, 25'd2019671, -25'd3168111, -25'd2376083, -25'd4197747, -25'd2455286, -25'd356412, -25'd3247314}, '{25'd1980069, 25'd2455286, -25'd1742461, -25'd2692894, 25'd3445321, 25'd1504853, -25'd3960139, -25'd2772097, 25'd2296881}, '{-25'd4237349, 25'd4039342, 25'd3128510, -25'd3722530, -25'd1940468, 25'd4593761, 25'd3999740, 25'd752426, -25'd1861265}, '{-25'd2296881, 25'd1267244, -25'd2296881, 25'd4831369, -25'd4316551, 25'd1504853, 25'd4593761, -25'd4474957, 25'd2336482}, '{-25'd2811699, 25'd3762132, -25'd4435355, 25'd1782062, -25'd2217678, -25'd3326517, 25'd1742461, 25'd118804, 25'd3405719}, '{-25'd5029376, 25'd2415685, -25'd752426, 25'd1821664, -25'd1346447, 25'd1029636, 25'd4237349, 25'd3286915, 25'd3524524}}, '{'{-25'd475217, 25'd4276950, 25'd3999740, -25'd3722530, 25'd1148440, -25'd4752167, -25'd1029636, -25'd3564125, 25'd4712565}, '{25'd0, 25'd3920537, -25'd1742461, 25'd3286915, -25'd2059272, 25'd1346447, 25'd3247314, -25'd1544454, -25'd2257279}, '{-25'd2772097, -25'd1663258, 25'd2772097, 25'd950433, -25'd2296881, 25'd554419, -25'd4316551, -25'd2534489, 25'd3920537}, '{25'd1227643, 25'd1148440, 25'd1504853, -25'd3326517, 25'd1069237, -25'd2296881, 25'd356412, -25'd1386049, 25'd435615}, '{25'd2653293, -25'd3207712, -25'd4276950, 25'd39601, 25'd3564125, -25'd3880936, 25'd514818, 25'd4474957, 25'd3841335}, '{-25'd3920537, -25'd4633362, -25'd1346447, 25'd475217, -25'd1544454, 25'd4672964, 25'd3643328, 25'd2613692, -25'd792028}, '{-25'd1623657, -25'd712825, -25'd1702860, -25'd2098874, 25'd475217, -25'd4316551, -25'd752426, -25'd4712565, -25'd3643328}, '{25'd910832, 25'd3999740, -25'd4197747, -25'd3484922, 25'd1900867, 25'd4356153, 25'd2811699, 25'd4593761, -25'd4276950}, '{25'd2851300, 25'd2178076, -25'd792028, -25'd118804, 25'd1900867, 25'd2376083, 25'd1108839, 25'd1425650, -25'd3207712}}},
    '{'{'{25'd3734212, 25'd1806877, 25'd1847030, 25'd2248558, -25'd3453142, -25'd1445501, 25'd2449322, 25'd3212225, 25'd4256199}, '{-25'd4617574, 25'd1405349, -25'd4175893, 25'd682598, 25'd4537268, 25'd722751, 25'd2248558, -25'd3453142, 25'd1847030}, '{25'd762904, -25'd2810697, 25'd4577421, -25'd2288711, 25'd1726571, 25'd3533448, -25'd2087946, -25'd401528, 25'd3774365}, '{-25'd1164432, 25'd2128099, 25'd2288711, 25'd441681, -25'd3734212, 25'd4256199, 25'd40153, -25'd401528, -25'd2850850}, '{25'd2971308, -25'd2168252, -25'd2007641, -25'd2489475, 25'd2208405, 25'd5099408, -25'd1405349, -25'd602292, 25'd2369016}, '{-25'd2087946, -25'd3854670, -25'd1164432, 25'd4778185, 25'd4015282, 25'd2168252, 25'd4697880, -25'd3131920, 25'd3894823}, '{25'd4978949, 25'd2128099, -25'd2409169, 25'd1043973, 25'd4898644, 25'd1124279, 25'd3212225, -25'd3774365, 25'd4778185}, '{-25'd160611, -25'd2047794, 25'd1405349, 25'd3091767, 25'd4336504, -25'd562139, 25'd602292, -25'd4456963, 25'd3011461}, '{-25'd4055434, -25'd923515, 25'd3814518, 25'd883362, -25'd1646265, -25'd3573601, -25'd963668, 25'd1806877, 25'd3372837}}, '{'{25'd2128099, 25'd843209, -25'd3292531, 25'd2168252, 25'd4135740, 25'd120458, -25'd4697880, -25'd4537268, 25'd722751}, '{-25'd2489475, -25'd3814518, -25'd843209, -25'd1806877, 25'd2690239, -25'd40153, 25'd3172072, 25'd4617574, 25'd481834}, '{-25'd1726571, 25'd3131920, -25'd1766724, -25'd4175893, 25'd120458, -25'd1325043, 25'd1806877, -25'd1686418, 25'd4336504}, '{-25'd2168252, 25'd843209, -25'd2128099, -25'd1084126, 25'd4497115, 25'd2609933, 25'd1325043, 25'd1847030, -25'd1606113}, '{25'd1325043, -25'd1606113, 25'd521987, 25'd2409169, 25'd4015282, 25'd1325043, -25'd441681, 25'd4296351, -25'd1284890}, '{-25'd2449322, 25'd3131920, -25'd3533448, 25'd3894823, 25'd4537268, 25'd3493295, 25'd1325043, -25'd3934976, 25'd3774365}, '{25'd4738032, -25'd441681, 25'd4577421, -25'd2810697, 25'd3292531, -25'd2569780, -25'd4336504, -25'd3533448, 25'd3212225}, '{-25'd1686418, 25'd80306, -25'd3734212, 25'd2087946, 25'd2128099, 25'd2850850, 25'd602292, 25'd3734212, 25'd1043973}, '{-25'd1847030, -25'd1525807, 25'd40153, 25'd2931156, -25'd1204584, -25'd883362, 25'd2891003, -25'd2810697, -25'd4095587}}, '{'{25'd1967488, 25'd2168252, -25'd3372837, -25'd200764, -25'd2810697, 25'd1847030, 25'd3854670, -25'd120458, 25'd3814518}, '{-25'd1124279, -25'd4456963, 25'd3172072, 25'd80306, -25'd2409169, 25'd0, 25'd4216046, 25'd1244737, 25'd2168252}, '{-25'd4095587, 25'd3131920, 25'd1043973, -25'd1204584, 25'd4216046, -25'd321223, -25'd2609933, -25'd602292, -25'd4898644}, '{25'd602292, -25'd4015282, 25'd562139, -25'd3854670, -25'd2369016, 25'd4818338, -25'd4818338, 25'd481834, 25'd883362}, '{-25'd3493295, 25'd4015282, 25'd4376657, -25'd2369016, 25'd1405349, -25'd2409169, 25'd3131920, -25'd1043973, -25'd3493295}, '{25'd2369016, 25'd4697880, 25'd0, -25'd2931156, -25'd1164432, 25'd3894823, -25'd562139, 25'd1284890, 25'd40153}, '{-25'd4135740, -25'd1606113, 25'd4657727, 25'd2891003, -25'd4216046, 25'd120458, 25'd4216046, -25'd3774365, -25'd4898644}, '{-25'd2609933, -25'd2690239, -25'd3854670, 25'd1043973, 25'd4256199, 25'd2971308, 25'd3573601, 25'd2931156, 25'd4738032}, '{-25'd2770544, -25'd1847030, -25'd4738032, -25'd3372837, -25'd4416810, 25'd1124279, -25'd4416810, -25'd2489475, -25'd3894823}}},
    '{'{'{-25'd3568488, 25'd3487386, -25'd729918, -25'd3284631, 25'd567714, 25'd1419285, 25'd3365733, -25'd364959, 25'd3487386}, '{-25'd3081876, -25'd1257081, -25'd3811794, 25'd4257855, 25'd4460610, -25'd2716917, 25'd4947222, 25'd2311407, -25'd81102}, '{-25'd1946448, -25'd405510, -25'd3527937, -25'd1865346, -25'd364959, 25'd527163, -25'd851571, -25'd1905897, 25'd3162978}, '{25'd932673, 25'd811020, 25'd2351958, -25'd2068101, -25'd4257855, 25'd2149203, -25'd3406284, -25'd608265, -25'd4379508}, '{-25'd3730692, 25'd729918, -25'd4298406, 25'd3203529, -25'd1946448, 25'd3081876, -25'd1257081, 25'd4298406, -25'd1419285}, '{25'd3568488, 25'd3325182, -25'd1297632, 25'd3365733, -25'd3122427, 25'd3203529, 25'd81102, 25'd446061, 25'd2879121}, '{-25'd1216530, 25'd1743693, -25'd4703916, 25'd567714, -25'd1135428, 25'd2270856, 25'd4744467, 25'd3527937, -25'd2311407}, '{25'd932673, 25'd4582263, -25'd1175979, -25'd486612, -25'd2392509, 25'd364959, -25'd2838570, 25'd1459836, 25'd3041325}, '{-25'd3162978, 25'd364959, 25'd283857, 25'd405510, -25'd3811794, 25'd364959, 25'd4703916, 25'd2838570, 25'd3203529}}, '{'{25'd4947222, -25'd3568488, 25'd364959, 25'd3730692, 25'd4866120, 25'd1905897, -25'd3527937, -25'd932673, 25'd4014549}, '{25'd3406284, 25'd648816, -25'd1622040, -25'd2514162, 25'd2189754, 25'd364959, 25'd2433060, -25'd1135428, -25'd2473611}, '{25'd1419285, -25'd3649590, -25'd1013775, 25'd2230305, 25'd324408, 25'd1905897, 25'd932673, 25'd811020, -25'd2635815}, '{25'd4420059, -25'd1257081, -25'd2068101, 25'd2798019, -25'd2068101, 25'd2716917, 25'd2757468, 25'd1946448, 25'd2514162}, '{25'd2473611, 25'd1824795, -25'd81102, -25'd4338957, 25'd405510, -25'd2514162, 25'd4136202, 25'd3730692, -25'd2960223}, '{-25'd2716917, -25'd2716917, -25'd2838570, 25'd5149977, 25'd2595264, 25'd608265, -25'd405510, 25'd4582263, 25'd3325182}, '{25'd4136202, 25'd4866120, 25'd202755, 25'd0, 25'd4501161, -25'd2514162, -25'd3852345, 25'd3609039, -25'd4420059}, '{25'd2798019, 25'd1865346, -25'd4541712, 25'd811020, 25'd4420059, 25'd527163, -25'd1216530, -25'd2514162, -25'd1581489}, '{25'd3649590, 25'd1824795, -25'd729918, 25'd3527937, -25'd1946448, 25'd1419285, 25'd1175979, -25'd3122427, -25'd1703142}}, '{'{-25'd4460610, 25'd1459836, -25'd3609039, 25'd202755, -25'd608265, 25'd4257855, -25'd1662591, -25'd2757468, -25'd1054326}, '{25'd4257855, -25'd3203529, -25'd4257855, -25'd3649590, 25'd4744467, 25'd40551, -25'd1338183, 25'd973224, -25'd4866120}, '{-25'd2757468, -25'd1703142, -25'd2554713, 25'd3122427, -25'd2189754, 25'd3852345, 25'd1703142, 25'd1905897, -25'd3730692}, '{-25'd1419285, -25'd4460610, 25'd4095651, 25'd2798019, -25'd2270856, 25'd4541712, 25'd1338183, -25'd4501161, -25'd364959}, '{-25'd3487386, 25'd324408, -25'd1865346, -25'd2757468, -25'd283857, 25'd1581489, 25'd4257855, 25'd1135428, -25'd4703916}, '{25'd4906671, 25'd2798019, 25'd3446835, -25'd3933447, -25'd243306, 25'd3081876, 25'd1378734, -25'd2311407, 25'd1703142}, '{25'd0, -25'd1622040, 25'd3365733, 25'd4663365, 25'd1622040, 25'd1865346, 25'd2149203, -25'd3365733, 25'd811020}, '{25'd2595264, 25'd0, -25'd1297632, 25'd3244080, -25'd4785018, 25'd2392509, -25'd2514162, -25'd121653, -25'd446061}, '{-25'd324408, -25'd1459836, 25'd3446835, 25'd3325182, 25'd2108652, -25'd446061, 25'd648816, -25'd4541712, -25'd4338957}}},
    '{'{'{25'd1013206, -25'd932149, 25'd1864299, 25'd1540073, 25'd3242258, -25'd2796448, -25'd2391166, 25'd1702186, -25'd3242258}, '{-25'd4214936, 25'd2958561, -25'd1702186, -25'd4498634, 25'd2836976, -25'd3039617, -25'd3485428, 25'd2310109, 25'd1337432}, '{-25'd2229053, -25'd4052823, -25'd4458105, 25'd3323315, 25'd3931238, 25'd1661657, 25'd1499545, -25'd283698, 25'd4255464}, '{-25'd486339, 25'd1783242, 25'd243169, -25'd4377049, -25'd729508, -25'd4701275, 25'd4174408, -25'd2715391, -25'd2715391}, '{25'd1783242, 25'd4093351, 25'd1256375, 25'd2147996, 25'd1377960, -25'd2147996, -25'd3525956, -25'd3647541, -25'd1580601}, '{-25'd1215847, -25'd2147996, -25'd688980, 25'd3931238, 25'd1459016, -25'd1296903, -25'd4660747, -25'd2715391, 25'd1864299}, '{25'd1459016, 25'd2269581, -25'd2553279, 25'd4012295, 25'd364754, 25'd3688069, -25'd3971767, 25'd2877504, -25'd1823770}, '{25'd2755920, 25'd2715391, -25'd3444900, -25'd2107468, 25'd4336521, -25'd1945355, 25'd526867, 25'd1945355, 25'd1256375}, '{25'd2634335, -25'd891621, -25'd1256375, 25'd1783242, -25'd4174408, 25'd2796448, -25'd2147996, -25'd3323315, 25'd2755920}}, '{'{-25'd3080146, -25'd1945355, -25'd3120674, 25'd4417577, -25'd2593807, -25'd405282, -25'd1742714, -25'd1702186, 25'd486339}, '{-25'd2269581, 25'd324226, 25'd891621, -25'd3525956, 25'd3769125, -25'd2431694, -25'd1864299, 25'd2026412, -25'd2674863}, '{-25'd1134790, 25'd3890710, 25'd2918033, 25'd3282787, 25'd1256375, 25'd729508, -25'd4863388, -25'd40528, 25'd1418488}, '{25'd3242258, 25'd2755920, -25'd2999089, -25'd2107468, 25'd526867, -25'd5187614, 25'd81056, -25'd2593807, -25'd324226}, '{-25'd1013206, 25'd3323315, -25'd3323315, -25'd3850182, 25'd4741803, -25'd4133880, -25'd3769125, 25'd2391166, -25'd1621129}, '{25'd3809654, -25'd3080146, 25'd4822859, -25'd2512750, -25'd1621129, -25'd4255464, 25'd4174408, -25'd2107468, 25'd4255464}, '{25'd1459016, -25'd3282787, 25'd486339, 25'd4944444, 25'd688980, -25'd5147085, 25'd1418488, -25'd1377960, -25'd729508}, '{-25'd1134790, -25'd4174408, -25'd1134790, -25'd2107468, 25'd2107468, -25'd486339, -25'd4701275, -25'd2391166, 25'd688980}, '{-25'd2553279, 25'd3809654, 25'd607923, 25'd2553279, -25'd4052823, -25'd4620218, -25'd243169, 25'd2836976, 25'd81056}}, '{'{25'd4944444, -25'd202641, -25'd2026412, 25'd81056, -25'd1499545, -25'd1459016, 25'd1621129, -25'd4741803, -25'd1134790}, '{-25'd202641, 25'd3161202, -25'd3809654, 25'd851093, -25'd1621129, 25'd891621, 25'd162113, 25'd2229053, 25'd3688069}, '{25'd2472222, 25'd4741803, 25'd729508, -25'd4377049, -25'd770036, -25'd2269581, -25'd202641, -25'd1580601, -25'd1256375}, '{-25'd2472222, -25'd81056, 25'd1985883, 25'd2310109, -25'd4295992, -25'd4822859, -25'd2958561, 25'd4539162, 25'd3161202}, '{25'd688980, 25'd2431694, -25'd932149, 25'd2310109, 25'd5147085, -25'd4498634, 25'd3525956, 25'd1904827, 25'd3890710}, '{25'd2715391, 25'd3769125, -25'd2593807, 25'd2796448, 25'd5147085, 25'd3120674, 25'd1945355, -25'd3080146, -25'd3242258}, '{-25'd1418488, 25'd2431694, -25'd4417577, -25'd2350637, -25'd2066940, 25'd3485428, 25'd3080146, -25'd5187614, 25'd2391166}, '{-25'd162113, -25'd2269581, 25'd4903916, 25'd729508, 25'd2674863, -25'd729508, 25'd648452, -25'd4052823, -25'd2836976}, '{-25'd1459016, -25'd1580601, 25'd2188524, -25'd567395, 25'd3728597, -25'd3323315, -25'd972678, 25'd162113, -25'd2674863}}},
    '{'{'{-25'd2555604, 25'd3132676, 25'd1442680, -25'd700730, 25'd1731216, 25'd1360241, 25'd3009018, 25'd1071705, -25'd2390727}, '{25'd1154144, 25'd0, 25'd2596824, 25'd4863892, -25'd2102191, 25'd1566338, 25'd2679263, -25'd370975, -25'd2473165}, '{-25'd3915845, -25'd1401460, 25'd1360241, 25'd4575356, 25'd2761701, 25'd659511, 25'd2555604, -25'd2514385, 25'd5069989}, '{-25'd4946331, -25'd948047, 25'd1071705, 25'd659511, -25'd3462432, 25'd3750968, -25'd3998284, -25'd4534137, 25'd4781453}, '{25'd3173896, -25'd2349507, -25'd2267068, 25'd3750968, -25'd3792187, -25'd4369259, -25'd4369259, -25'd2844140, -25'd1195363}, '{25'd2885360, 25'd2761701, -25'd370975, 25'd4410478, -25'd3462432, 25'd4163162, -25'd3173896, -25'd4410478, 25'd659511}, '{25'd3009018, -25'd2720482, 25'd1360241, 25'd3215115, 25'd3050237, -25'd3256335, 25'd123658, 25'd2967799, -25'd412194}, '{-25'd824388, -25'd3792187, -25'd4740234, -25'd3379993, 25'd4987550, -25'd453414, 25'd2184630, 25'd3421212, -25'd2390727}, '{25'd1648777, -25'd3091457, -25'd906827, 25'd1071705, -25'd247317, 25'd1854874, -25'd247317, -25'd3957065, -25'd2638043}}, '{'{-25'd4328040, 25'd453414, -25'd4863892, 25'd4204381, 25'd4080723, 25'd4863892, -25'd4699014, 25'd2514385, 25'd2431946}, '{25'd3338773, 25'd2679263, -25'd989266, 25'd1689996, 25'd3627309, -25'd1689996, -25'd659511, -25'd3256335, 25'd1648777}, '{-25'd3915845, -25'd494633, 25'd2720482, -25'd4245601, -25'd2225849, 25'd494633, 25'd3009018, -25'd3668529, 25'd577072}, '{-25'd3998284, 25'd577072, 25'd535853, 25'd4410478, 25'd4657795, -25'd824388, -25'd41219, 25'd2885360, -25'd82439}, '{25'd3215115, -25'd3998284, -25'd2349507, -25'd1195363, -25'd2885360, -25'd1442680, 25'd3421212, -25'd2390727, -25'd41219}, '{25'd1607558, -25'd1854874, -25'd1937313, 25'd41219, -25'd288536, 25'd41219, -25'd865608, 25'd206097, -25'd4451698}, '{-25'd1731216, 25'd4039504, -25'd4616576, -25'd4369259, 25'd865608, 25'd3173896, -25'd82439, -25'd3379993, -25'd4328040}, '{25'd2060971, -25'd1896094, -25'd164878, -25'd1277802, -25'd412194, -25'd1360241, 25'd3750968, 25'd3544871, 25'd5028770}, '{-25'd2638043, 25'd3503651, -25'd1525119, 25'd741950, 25'd5234867, 25'd1360241, 25'd3462432, -25'd2844140, 25'd3792187}}, '{'{-25'd2802921, -25'd1442680, -25'd5111209, -25'd1030486, 25'd1112924, 25'd1978532, -25'd2431946, -25'd3050237, -25'd2473165}, '{-25'd1566338, -25'd1648777, 25'd4492917, 25'd1689996, 25'd1772435, -25'd494633, -25'd453414, 25'd1030486, -25'd164878}, '{25'd1937313, 25'd41219, -25'd906827, 25'd4451698, 25'd3503651, 25'd3750968, 25'd2885360, -25'd3462432, -25'd1731216}, '{-25'd1401460, 25'd329755, 25'd2802921, 25'd4410478, -25'd4575356, -25'd1195363, 25'd288536, -25'd1319022, 25'd288536}, '{-25'd4163162, -25'd4822673, 25'd3132676, -25'd2926579, -25'd2143410, 25'd1689996, -25'd206097, -25'd2638043, 25'd3998284}, '{25'd4039504, -25'd4410478, -25'd3379993, -25'd3050237, 25'd370975, 25'd3009018, -25'd1854874, 25'd2349507, -25'd3833406}, '{-25'd3709748, -25'd2679263, 25'd1937313, -25'd3215115, -25'd1401460, 25'd370975, 25'd2225849, 25'd206097, -25'd1236583}, '{25'd123658, -25'd2596824, 25'd1896094, 25'd2638043, -25'd1154144, 25'd4369259, -25'd1566338, 25'd1401460, -25'd3091457}, '{25'd4863892, 25'd247317, 25'd3998284, -25'd2679263, -25'd2638043, 25'd2019752, 25'd3627309, 25'd4080723, 25'd2225849}}},
    '{'{'{25'd4037190, 25'd2580472, 25'd1331856, 25'd3496123, 25'd4786359, 25'd1706441, -25'd2455610, -25'd4744738, -25'd83241}, '{25'd2580472, -25'd1539959, 25'd541067, -25'd2164267, -25'd832410, -25'd4411774, 25'd3038297, -25'd166482, -25'd1206995}, '{-25'd4245292, -25'd124862, 25'd2663713, 25'd3204779, -25'd3246400, -25'd2996677, 25'd4078810, 25'd4703118, 25'd582687}, '{-25'd3537744, 25'd4411774, 25'd4619877, 25'd3038297, 25'd624308, 25'd332964, -25'd832410, 25'd3371261, -25'd2081026}, '{25'd1082133, -25'd3870708, -25'd1456718, -25'd2830195, -25'd2705333, 25'd5202564, -25'd2497231, 25'd5119323, 25'd1623200}, '{-25'd4453395, 25'd1623200, -25'd1123754, 25'd4370154, 25'd1165374, -25'd3787467, 25'd665928, 25'd3745846, 25'd707549}, '{-25'd4370154, 25'd2788574, 25'd1415097, -25'd4536636, -25'd2039405, 25'd1082133, -25'd1123754, 25'd582687, -25'd499446}, '{-25'd2413990, -25'd2081026, 25'd2497231, 25'd1706441, -25'd2996677, 25'd374585, 25'd3371261, 25'd1373477, 25'd3537744}, '{25'd915651, -25'd1165374, 25'd2330749, 25'd2289128, 25'd3204779, 25'd332964, -25'd1123754, 25'd1373477, -25'd2372369}}, '{'{-25'd3288020, -25'd2705333, -25'd4453395, 25'd665928, 25'd4370154, -25'd4495015, 25'd1082133, -25'd2455610, -25'd2205887}, '{25'd4411774, -25'd2913436, -25'd1206995, -25'd2788574, -25'd3204779, -25'd2913436, -25'd790790, -25'd957272, 25'd1290236}, '{-25'd208103, 25'd4744738, -25'd2413990, 25'd3745846, 25'd3246400, -25'd3995569, -25'd2913436, 25'd4578256, -25'd4786359}, '{25'd1748062, -25'd3329641, -25'd2413990, 25'd665928, -25'd3995569, -25'd1123754, -25'd249723, -25'd2871815, -25'd4037190}, '{-25'd3995569, 25'd4578256, 25'd4578256, 25'd4619877, 25'd2663713, 25'd5285805, -25'd3412882, 25'd4703118, -25'd2372369}, '{25'd3121538, 25'd4661497, 25'd3079918, -25'd3662605, 25'd915651, -25'd582687, 25'd41621, -25'd2746954, 25'd499446}, '{25'd4578256, 25'd998892, -25'd1623200, -25'd1872923, 25'd1706441, 25'd4245292, -25'd1664820, 25'd2497231, -25'd4536636}, '{25'd208103, -25'd1748062, 25'd2746954, -25'd2039405, -25'd1706441, 25'd4245292, -25'd790790, 25'd5077702, 25'd2580472}, '{-25'd624308, 25'd83241, 25'd4411774, -25'd3288020, -25'd2413990, 25'd4827979, 25'd3579364, -25'd541067, -25'd2871815}}, '{'{25'd2497231, -25'd2330749, 25'd4370154, -25'd2247508, 25'd208103, -25'd4453395, -25'd1373477, -25'd2497231, 25'd3870708}, '{25'd1165374, 25'd1706441, 25'd4495015, 25'd4578256, 25'd2039405, 25'd1706441, -25'd4536636, 25'd832410, 25'd332964}, '{25'd1914544, 25'd3163159, 25'd3496123, -25'd4078810, 25'd4453395, -25'd1872923, 25'd3912328, -25'd790790, -25'd4411774}, '{-25'd208103, 25'd4536636, 25'd1290236, -25'd1498338, 25'd4453395, 25'd499446, -25'd2871815, 25'd3454503, 25'd2746954}, '{-25'd1664820, 25'd3371261, 25'd4162051, 25'd1748062, -25'd1082133, 25'd2705333, 25'd166482, 25'd249723, -25'd2538851}, '{-25'd4786359, -25'd4286913, 25'd374585, -25'd3371261, 25'd957272, 25'd374585, 25'd2622092, -25'd4245292, 25'd3121538}, '{25'd2622092, -25'd1123754, -25'd4370154, 25'd4370154, 25'd2871815, 25'd957272, -25'd874031, 25'd1373477, -25'd41621}, '{25'd2372369, -25'd2122646, 25'd4286913, 25'd249723, 25'd3121538, -25'd2788574, 25'd4619877, -25'd998892, -25'd249723}, '{25'd3745846, -25'd2247508, -25'd457826, 25'd3038297, -25'd4078810, -25'd541067, -25'd4453395, 25'd3204779, 25'd1831303}}},
    '{'{'{25'd2569086, 25'd4415617, 25'd3251500, 25'd2569086, -25'd2328234, -25'd1244401, -25'd762697, 25'd1404969, -25'd441562}, '{25'd1605679, 25'd4857178, 25'd1364827, -25'd1685963, 25'd441562, -25'd3893771, 25'd1003549, -25'd3090932, -25'd1525395}, '{25'd4616327, 25'd1284543, 25'd200710, 25'd2528944, 25'd3974055, 25'd1726105, -25'd802839, -25'd2569086, -25'd4335333}, '{-25'd3572635, -25'd4174765, -25'd2769796, -25'd2970506, 25'd3171216, -25'd642272, -25'd762697, 25'd2368376, -25'd1445111}, '{25'd3131074, 25'd1043691, -25'd3090932, -25'd2890222, -25'd3211358, -25'd1886673, 25'd682413, 25'd4656469, -25'd2809938}, '{25'd1966957, 25'd2328234, 25'd1364827, -25'd842981, 25'd2649370, -25'd2408518, -25'd1324685, 25'd4174765, -25'd3131074}, '{-25'd3010648, 25'd4495901, -25'd2809938, -25'd4857178, -25'd4776894, 25'd1485253, -25'd200710, 25'd963407, -25'd200710}, '{-25'd1485253, 25'd1445111, -25'd923265, 25'd842981, 25'd1404969, -25'd3612777, 25'd361278, -25'd4696611, 25'd4214907}, '{25'd3492351, 25'd4134623, 25'd1886673, -25'd2609228, -25'd4415617, 25'd4375475, -25'd200710, 25'd3612777, 25'd3693061}}, '{'{-25'd2528944, 25'd2769796, -25'd923265, -25'd2047240, -25'd2488802, -25'd3974055, 25'd2528944, 25'd4616327, 25'd1605679}, '{25'd682413, 25'd2007099, 25'd4214907, -25'd1404969, 25'd1204259, -25'd1806389, 25'd2609228, 25'd4696611, -25'd1525395}, '{25'd1003549, -25'd2127524, 25'd3131074, -25'd682413, 25'd1926815, 25'd2167666, 25'd2729654, -25'd2890222, -25'd2609228}, '{25'd4255049, 25'd4576185, 25'd3452209, -25'd441562, 25'd3652919, 25'd1123975, 25'd4335333, -25'd1083833, 25'd4335333}, '{25'd2007099, -25'd3733203, -25'd1685963, 25'd1083833, 25'd1284543, 25'd1083833, 25'd3933913, 25'd3452209, -25'd401420}, '{25'd2127524, 25'd2930364, 25'd2127524, -25'd3452209, -25'd3412067, -25'd3893771, -25'd642272, -25'd4014197, 25'd1284543}, '{-25'd3251500, -25'd1364827, 25'd963407, 25'd1364827, -25'd3532493, 25'd4656469, 25'd200710, 25'd802839, 25'd1485253}, '{-25'd2769796, 25'd3131074, 25'd2408518, 25'd2729654, 25'd1445111, 25'd1364827, 25'd4335333, -25'd602130, -25'd3733203}, '{-25'd1244401, 25'd4335333, 25'd1083833, 25'd5017746, -25'd4455759, 25'd2007099, 25'd2448660, 25'd963407, 25'd200710}}, '{'{25'd3532493, -25'd4134623, -25'd4455759, 25'd5017746, -25'd3452209, 25'd2809938, -25'd2769796, -25'd240852, -25'd3773345}, '{25'd401420, 25'd2047240, 25'd2368376, 25'd3452209, 25'd2007099, 25'd2207808, 25'd3291642, -25'd3974055, -25'd4817036}, '{-25'd2649370, -25'd682413, -25'd1926815, -25'd1766247, -25'd3572635, 25'd200710, 25'd1645821, 25'd4054339, 25'd602130}, '{-25'd2288092, 25'd2368376, 25'd2769796, -25'd561988, -25'd4054339, 25'd1565537, -25'd1204259, 25'd4495901, 25'd1605679}, '{25'd280994, -25'd4214907, -25'd682413, 25'd3572635, 25'd1244401, 25'd3251500, 25'd4214907, 25'd1485253, -25'd1324685}, '{25'd3131074, -25'd401420, -25'd1324685, 25'd1445111, -25'd2047240, 25'd4536043, 25'd481704, -25'd1886673, -25'd762697}, '{25'd2087382, 25'd1685963, -25'd280994, 25'd4134623, -25'd2328234, -25'd2087382, -25'd3331784, -25'd1485253, -25'd3933913}, '{25'd1204259, -25'd1926815, 25'd1083833, -25'd1525395, -25'd883123, -25'd4576185, -25'd3010648, -25'd1485253, 25'd5098030}, '{25'd1685963, 25'd120426, 25'd4576185, 25'd2167666, 25'd4174765, 25'd441562, 25'd3612777, -25'd1726105, 25'd4656469}}},
    '{'{'{-25'd4009542, 25'd4358198, -25'd4881182, 25'd2266263, 25'd5404165, -25'd232437, 25'd755421, 25'd3718996, 25'd290547}, '{-25'd2963575, -25'd4648745, -25'd4300089, -25'd290547, -25'd581093, -25'd290547, -25'd3196012, 25'd1220295, -25'd3196012}, '{25'd2440591, -25'd2091935, 25'd2440591, -25'd1394623, 25'd5810931, -25'd581093, -25'd1104077, -25'd116219, -25'd2556809}, '{25'd2963575, 25'd3951433, 25'd4067651, 25'd697312, 25'd232437, 25'd1104077, 25'd2150044, -25'd3951433, 25'd3718996}, '{25'd4241979, 25'd2324372, 25'd4067651, 25'd7263663, -25'd813530, 25'd1917607, -25'd464874, 25'd2440591, -25'd3893324}, '{25'd3544668, -25'd2440591, -25'd581093, 25'd4823072, 25'd4358198, 25'd7379882, 25'd232437, 25'd3544668, 25'd3718996}, '{-25'd522984, -25'd581093, -25'd4939291, -25'd1801388, 25'd1278405, 25'd4067651, -25'd2324372, -25'd4706854, -25'd1394623}, '{-25'd2033826, -25'd1394623, -25'd4706854, 25'd2905465, -25'd3254121, 25'd3254121, 25'd1336514, -25'd290547, -25'd4358198}, '{25'd348656, -25'd4823072, -25'd2963575, -25'd2266263, -25'd1743279, 25'd2266263, -25'd3021684, 25'd987858, 25'd2731137}}, '{'{25'd3137903, 25'd4067651, -25'd871640, 25'd3312230, -25'd2556809, -25'd290547, -25'd232437, -25'd3312230, 25'd4532526}, '{-25'd1801388, 25'd4939291, -25'd2440591, 25'd5636603, 25'd755421, -25'd58109, 25'd4648745, 25'd2266263, -25'd116219}, '{-25'd3196012, -25'd1975716, -25'd2033826, -25'd290547, 25'd1743279, 25'd2905465, 25'd1104077, 25'd58109, -25'd2673028}, '{-25'd3486558, 25'd116219, 25'd232437, 25'd7089335, 25'd5520384, -25'd1568951, 25'd5927149, 25'd5636603, 25'd1394623}, '{-25'd1220295, 25'd2440591, 25'd3602777, 25'd58109, -25'd58109, 25'd4881182, 25'd348656, 25'd755421, 25'd4706854}, '{-25'd2150044, 25'd639202, -25'd1278405, 25'd174328, 25'd4300089, 25'd1220295, 25'd5694712, -25'd464874, -25'd2498700}, '{-25'd2440591, -25'd5927149, -25'd4939291, 25'd1801388, -25'd639202, -25'd3312230, 25'd3312230, 25'd2091935, 25'd639202}, '{-25'd755421, -25'd6043368, -25'd6217696, -25'd3951433, -25'd3951433, 25'd639202, -25'd2614919, -25'd2150044, -25'd2673028}, '{-25'd1104077, -25'd6682570, -25'd639202, -25'd3835214, -25'd522984, -25'd4881182, 25'd3777105, -25'd116219, -25'd4939291}}, '{'{25'd2731137, 25'd1510842, -25'd871640, 25'd2150044, 25'd5113619, 25'd2614919, -25'd1452733, -25'd2382482, -25'd697312}, '{25'd1975716, 25'd4300089, 25'd3196012, 25'd1917607, -25'd522984, -25'd1685170, 25'd871640, -25'd4532526, 25'd1975716}, '{25'd1568951, -25'd1685170, 25'd3777105, -25'd1336514, 25'd4823072, -25'd929749, -25'd522984, -25'd4241979, -25'd522984}, '{-25'd5055510, 25'd4416307, -25'd755421, 25'd6973117, 25'd5927149, 25'd1394623, 25'd0, 25'd4474417, 25'd3021684}, '{-25'd3137903, 25'd2731137, -25'd3312230, 25'd7147445, 25'd1975716, 25'd4009542, 25'd5810931, 25'd1162186, -25'd1452733}, '{-25'd929749, 25'd4241979, -25'd1859498, 25'd6217696, 25'd639202, 25'd813530, 25'd5985259, -25'd232437, 25'd1859498}, '{-25'd4881182, -25'd5927149, 25'd1917607, 25'd5055510, -25'd232437, 25'd813530, 25'd2033826, -25'd3196012, -25'd1336514}, '{-25'd6217696, -25'd581093, -25'd4300089, 25'd232437, -25'd3312230, -25'd2498700, 25'd3893324, 25'd2614919, 25'd1278405}, '{-25'd2847356, -25'd3254121, 25'd58109, -25'd1685170, -25'd464874, -25'd639202, -25'd4183870, -25'd4125761, 25'd2382482}}},
    '{'{'{-25'd1366584, -25'd341646, -25'd3032108, -25'd3501871, 25'd597880, -25'd2647756, -25'd1708230, 25'd1281172, 25'd3074814}, '{-25'd2989402, -25'd3758106, -25'd768703, 25'd3160225, 25'd1964464, 25'd3886223, 25'd4355986, 25'd4057046, -25'd3373754}, '{-25'd1451995, 25'd2007170, 25'd4996572, -25'd1708230, 25'd1409290, 25'd2263405, 25'd2306110, -25'd2818579, 25'd4612221}, '{-25'd2135287, -25'd4057046, -25'd768703, 25'd42706, 25'd811409, 25'd2946696, 25'd4783044, -25'd1708230, 25'd4099752}, '{-25'd3245637, 25'd341646, -25'd1921759, 25'd3672694, 25'd1366584, 25'd1323878, 25'd0, -25'd4057046, -25'd768703}, '{25'd2775873, 25'd2434228, 25'd4014340, -25'd982232, 25'd4484103, -25'd3843517, -25'd4185163, -25'd4484103, 25'd1921759}, '{-25'd341646, -25'd1451995, -25'd4441398, -25'd1793641, -25'd3074814, -25'd4398692, -25'd298940, -25'd3032108, -25'd1238467}, '{-25'd2946696, 25'd4313280, -25'd2605051, 25'd2818579, -25'd982232, -25'd811409, -25'd4142457, -25'd3117519, 25'd1366584}, '{-25'd1366584, -25'd2946696, 25'd3160225, -25'd2861285, -25'd4014340, 25'd725998, 25'd4654926, -25'd640586, 25'd128117}}, '{'{25'd4185163, -25'd3928929, -25'd3245637, -25'd2775873, 25'd256234, 25'd170823, 25'd3758106, -25'd1494701, -25'd2391522}, '{25'd2775873, 25'd1921759, 25'd1793641, -25'd896821, -25'd4654926, 25'd4398692, 25'd256234, 25'd3544577, 25'd2220699}, '{-25'd1366584, 25'd4441398, -25'd2434228, 25'd3373754, -25'd1451995, -25'd4654926, 25'd3501871, 25'd4313280, 25'd4014340}, '{25'd3544577, 25'd384352, 25'd4142457, -25'd1921759, 25'd1580113, 25'd2434228, 25'd3629988, 25'd4526809, 25'd85411}, '{25'd4227869, -25'd512469, -25'd1921759, 25'd4057046, 25'd939526, -25'd3843517, -25'd3117519, -25'd3160225, 25'd2605051}, '{25'd640586, -25'd3928929, -25'd2989402, -25'd3288342, 25'd3758106, 25'd3459165, -25'd4612221, -25'd3160225, -25'd1750936}, '{25'd1110349, 25'd3672694, 25'd256234, 25'd4227869, 25'd4355986, -25'd4014340, -25'd768703, -25'd1366584, -25'd2135287}, '{-25'd3160225, 25'd3971634, -25'd1366584, 25'd2861285, 25'd213529, 25'd2733168, -25'd4654926, -25'd1665524, 25'd1836347}, '{25'd2733168, -25'd3373754, 25'd3160225, 25'd2135287, 25'd1195761, -25'd4313280, -25'd1879053, -25'd3672694, 25'd4526809}}, '{'{-25'd85411, 25'd3459165, 25'd4355986, -25'd1793641, 25'd2049876, -25'd1323878, 25'd3758106, -25'd1879053, 25'd4014340}, '{-25'd1281172, 25'd170823, -25'd2562345, 25'd170823, 25'd170823, -25'd3459165, 25'd2263405, -25'd1921759, 25'd1153055}, '{-25'd2049876, -25'd2733168, 25'd3843517, 25'd1067644, 25'd42706, 25'd4313280, -25'd3501871, -25'd683292, -25'd1793641}, '{-25'd2861285, 25'd1537407, 25'd4185163, 25'd768703, -25'd4142457, -25'd3245637, -25'd4057046, 25'd811409, -25'd1153055}, '{25'd4484103, 25'd683292, 25'd213529, -25'd1067644, -25'd213529, -25'd3459165, 25'd2647756, -25'd3245637, 25'd3928929}, '{25'd341646, -25'd2220699, 25'd1323878, 25'd5423630, -25'd4099752, 25'd0, 25'd3715400, -25'd3843517, 25'd4313280}, '{-25'd4484103, 25'd3416460, 25'd2135287, -25'd1281172, 25'd5081984, 25'd2135287, -25'd1494701, 25'd1793641, -25'd4014340}, '{25'd768703, 25'd4227869, -25'd85411, 25'd4868455, 25'd1708230, 25'd42706, 25'd1879053, 25'd213529, -25'd2903991}, '{25'd1879053, 25'd1750936, 25'd683292, 25'd3160225, 25'd2605051, 25'd3416460, 25'd2861285, 25'd256234, -25'd2135287}}},
    '{'{'{25'd3967836, -25'd2946413, -25'd1571420, -25'd1414278, -25'd78571, -25'd667854, 25'd1964275, 25'd3457124, -25'd3103555}, '{-25'd2985698, 25'd4635689, -25'd3299982, -25'd471426, -25'd1532135, 25'd3732123, -25'd4517833, 25'd2278559, 25'd2632129}, '{-25'd4399976, 25'd1374993, -25'd4871402, -25'd1571420, 25'd2278559, -25'd2278559, -25'd3535695, 25'd1649991, -25'd1807133}, '{-25'd3771408, 25'd3732123, 25'd4007121, 25'd4242834, 25'd3024984, -25'd3417839, 25'd4399976, 25'd4360691, -25'd1296422}, '{25'd1846419, -25'd4832117, 25'd2278559, 25'd117857, -25'd4832117, -25'd4046407, -25'd3417839, -25'd4557118, -25'd903567}, '{-25'd4635689, 25'd2749985, 25'd2317845, 25'd4557118, -25'd2671414, -25'd39286, 25'd1532135, 25'd471426, -25'd2749985}, '{-25'd471426, -25'd1807133, 25'd903567, -25'd1296422, 25'd2003561, 25'd2003561, 25'd3771408, 25'd1846419, 25'd4517833}, '{25'd4164263, 25'd117857, -25'd3103555, 25'd4124978, -25'd4124978, 25'd4242834, -25'd235713, 25'd1649991, -25'd942852}, '{25'd3260697, 25'd3535695, -25'd2907127, -25'd1767848, -25'd2946413, 25'd1099994, 25'd3692837, -25'd4871402, -25'd2592843}}, '{'{-25'd2396416, -25'd3221411, -25'd3574981, 25'd1099994, -25'd2514272, 25'd824996, -25'd3928550, 25'd3417839, 25'd3378553}, '{25'd2592843, 25'd2317845, -25'd1139280, -25'd353570, -25'd235713, -25'd2042846, -25'd4989259, 25'd1335707, 25'd2632129}, '{-25'd667854, 25'd3417839, 25'd3928550, 25'd785710, 25'd1767848, -25'd589283, -25'd2042846, -25'd235713, 25'd4557118}, '{-25'd785710, -25'd78571, -25'd4321405, -25'd3339268, -25'd3457124, -25'd4832117, 25'd3771408, 25'd3103555, -25'd392855}, '{-25'd1178565, 25'd1099994, 25'd274999, -25'd1296422, -25'd2199988, 25'd3103555, 25'd2828556, -25'd2592843, -25'd4871402}, '{-25'd549997, -25'd3378553, -25'd4478547, 25'd3221411, 25'd1296422, -25'd1610706, 25'd3574981, -25'd2710700, -25'd3496410}, '{25'd3574981, 25'd1453564, -25'd4164263, -25'd549997, 25'd1374993, -25'd471426, -25'd4282120, 25'd2003561, 25'd1689277}, '{25'd1532135, 25'd1414278, -25'd3574981, -25'd1728562, 25'd3928550, 25'd2514272, -25'd1492849, -25'd2435701, 25'd1492849}, '{25'd2199988, -25'd3810694, -25'd2632129, 25'd1335707, -25'd1021423, -25'd3221411, -25'd3024984, 25'd1689277, -25'd4871402}}, '{'{-25'd157142, -25'd2710700, 25'd3967836, -25'd1610706, -25'd4478547, -25'd471426, -25'd3732123, 25'd3535695, -25'd4753546}, '{-25'd3417839, -25'd2828556, -25'd4439262, -25'd1532135, 25'd510712, -25'd3299982, -25'd3299982, 25'd3928550, -25'd1414278}, '{25'd1649991, -25'd3103555, -25'd4792831, -25'd3810694, 25'd1335707, -25'd3967836, 25'd2592843, 25'd1964275, -25'd1099994}, '{-25'd1217851, -25'd4046407, -25'd746425, -25'd1846419, -25'd2789271, 25'd2632129, -25'd2671414, -25'd196428, -25'd3849979}, '{-25'd1217851, -25'd2985698, -25'd2867842, -25'd2160703, 25'd2435701, 25'd4596404, -25'd4989259, -25'd1571420, -25'd3260697}, '{-25'd2082132, -25'd3849979, 25'd3457124, -25'd4596404, 25'd1257136, 25'd2553558, 25'd510712, -25'd3339268, 25'd3103555}, '{-25'd3771408, 25'd864281, -25'd1532135, -25'd3299982, -25'd4046407, 25'd4321405, -25'd1649991, -25'd1492849, 25'd2985698}, '{-25'd2003561, 25'd3614266, 25'd3417839, 25'd3221411, 25'd3378553, 25'd1846419, 25'd2082132, -25'd2199988, -25'd2317845}, '{-25'd2946413, -25'd2514272, 25'd1060709, 25'd1532135, 25'd2592843, -25'd1767848, -25'd2632129, -25'd3614266, -25'd3260697}}},
    '{'{'{25'd2875092, -25'd498349, 25'd2453412, -25'd2185070, -25'd345011, 25'd4523478, 25'd4370140, 25'd4638482, 25'd4063464}, '{25'd2223405, 25'd4830155, 25'd1495048, -25'd728357, 25'd3373441, 25'd345011, -25'd3871791, 25'd3296772, -25'd1188371}, '{25'd3143434, -25'd2760088, -25'd2951761, 25'd4140133, 25'd805026, -25'd575018, -25'd4140133, -25'd191673, 25'd4255136}, '{-25'd1571717, -25'd3258438, 25'd1073368, 25'd3795122, 25'd3986794, 25'd766691, -25'd1495048, 25'd1801724, 25'd4140133}, '{-25'd1226706, 25'd2108401, 25'd4255136, 25'd268342, -25'd2645085, 25'd345011, 25'd4370140, -25'd2683419, 25'd2491747}, '{25'd3948460, -25'd881695, 25'd2760088, 25'd3335107, 25'd1380044, 25'd2645085, -25'd1840059, -25'd3526780, 25'd1226706}, '{-25'd4370140, -25'd1303375, 25'd3143434, -25'd1571717, 25'd3910125, -25'd1188371, 25'd3948460, 25'd4600147, 25'd1955063}, '{25'd4676817, 25'd1763390, 25'd76669, -25'd191673, 25'd230007, -25'd1188371, -25'd4063464, 25'd3411776, -25'd1226706}, '{-25'd3411776, -25'd3871791, -25'd498349, -25'd1878394, -25'd3028430, -25'd115004, 25'd2875092, 25'd3986794, 25'd1418379}}, '{'{25'd1725055, 25'd0, -25'd1878394, -25'd1111702, 25'd3450111, 25'd4063464, -25'd1725055, 25'd3220103, 25'd4025129}, '{-25'd1380044, 25'd498349, 25'd613353, -25'd2606750, -25'd4331806, -25'd2453412, 25'd153338, -25'd4293471, -25'd2606750}, '{-25'd2645085, -25'd3258438, -25'd1265041, 25'd4868489, 25'd3296772, 25'd3258438, -25'd1150037, -25'd1303375, 25'd306676}, '{25'd4600147, -25'd805026, 25'd4715151, 25'd613353, 25'd4370140, -25'd1456713, -25'd191673, -25'd1418379, -25'd3143434}, '{25'd3603449, 25'd881695, 25'd1341710, 25'd2875092, -25'd2031732, 25'd2070066, -25'd268342, 25'd3948460, -25'd3756787}, '{-25'd1341710, -25'd996699, -25'd1725055, -25'd1495048, 25'd2376743, 25'd3488445, 25'd2760088, -25'd4101798, 25'd2070066}, '{-25'd2951761, 25'd2836758, -25'd2415077, 25'd4063464, 25'd3105100, 25'd2606750, -25'd3488445, -25'd1725055, -25'd4753486}, '{25'd4025129, 25'd0, 25'd2108401, 25'd4370140, -25'd3028430, -25'd1111702, -25'd2185070, -25'd1303375, -25'd4676817}, '{-25'd3833456, 25'd3066765, 25'd1265041, 25'd3335107, 25'd2491747, 25'd1418379, 25'd3603449, -25'd1265041, 25'd4178467}}, '{'{25'd3450111, -25'd1533382, 25'd4446809, 25'd3718453, 25'd1993397, 25'd4600147, 25'd613353, 25'd2836758, 25'd0}, '{25'd2913427, 25'd2913427, 25'd191673, -25'd2683419, 25'd575018, -25'd766691, 25'd843360, -25'd115004, 25'd805026}, '{25'd2376743, 25'd1916728, -25'd843360, -25'd805026, 25'd2683419, 25'd2836758, 25'd1341710, -25'd1840059, -25'd2031732}, '{-25'd4830155, 25'd4523478, 25'd230007, 25'd4216802, 25'd3910125, -25'd1648386, -25'd153338, -25'd1916728, -25'd1303375}, '{25'd230007, 25'd2913427, 25'd4485144, 25'd881695, -25'd2990096, 25'd2031732, -25'd191673, 25'd306676, -25'd2453412}, '{-25'd1265041, 25'd1341710, 25'd2185070, -25'd958364, 25'd3641783, -25'd3871791, 25'd3526780, -25'd1955063, 25'd4101798}, '{-25'd4523478, 25'd4331806, -25'd2376743, -25'd115004, 25'd2721754, -25'd2108401, 25'd4178467, -25'd1801724, 25'd1840059}, '{25'd3258438, 25'd2530081, -25'd1456713, -25'd2108401, 25'd4178467, -25'd1763390, 25'd2261739, -25'd115004, -25'd4370140}, '{-25'd230007, 25'd2913427, 25'd345011, -25'd4025129, -25'd4331806, 25'd345011, 25'd2875092, 25'd1571717, -25'd2223405}}},
    '{'{'{-25'd4407048, -25'd440705, -25'd4186695, 25'd2864581, 25'd3158384, -25'd1248664, 25'd3378737, -25'd2130073, -25'd2644229}, '{-25'd146902, 25'd0, -25'd4260146, 25'd3966343, 25'd1836270, -25'd2644229, 25'd3819441, -25'd73451, -25'd3892892}, '{25'd3672540, 25'd3525638, -25'd514156, 25'd1028311, -25'd3452187, -25'd2717679, -25'd5288457, 25'd4260146, -25'd3305286}, '{25'd2130073, 25'd3084933, 25'd3892892, 25'd3452187, -25'd2644229, -25'd4480498, -25'd1028311, -25'd3378737, -25'd1395565}, '{-25'd3084933, 25'd3158384, 25'd2276975, -25'd587606, 25'd734508, -25'd734508, 25'd293803, -25'd1762819, -25'd4847752}, '{25'd3892892, -25'd4553949, 25'd4113244, -25'd4039794, -25'd73451, -25'd4407048, -25'd1469016, -25'd4113244, 25'd2130073}, '{-25'd7491981, -25'd2497327, -25'd6830924, -25'd6537121, -25'd2864581, -25'd4407048, -25'd8960997, -25'd5435359, -25'd9401702}, '{-25'd4333597, -25'd3084933, -25'd514156, -25'd7785784, -25'd8079587, -25'd3305286, -25'd3672540, -25'd6904375, -25'd1395565}, '{-25'd6243318, -25'd6977825, -25'd5582260, -25'd1689368, -25'd1689368, -25'd7785784, -25'd7418530, -25'd3084933, -25'd3158384}}, '{'{-25'd4627400, -25'd1028311, 25'd3599089, 25'd1395565, 25'd1469016, 25'd1762819, 25'd2130073, -25'd2350425, 25'd661057}, '{25'd0, 25'd3819441, 25'd3672540, 25'd2350425, 25'd4407048, 25'd3158384, 25'd4039794, -25'd3452187, 25'd1322114}, '{-25'd3819441, 25'd881410, -25'd293803, -25'd1689368, 25'd5435359, -25'd1542467, 25'd5215006, 25'd514156, 25'd734508}, '{-25'd2791130, 25'd3158384, 25'd146902, -25'd1615917, 25'd1689368, 25'd4039794, -25'd2056622, 25'd4333597, 25'd146902}, '{-25'd3452187, 25'd3011483, -25'd146902, 25'd73451, -25'd220352, 25'd514156, 25'd5141556, -25'd1101762, -25'd514156}, '{-25'd2130073, 25'd1322114, 25'd1028311, -25'd2497327, 25'd6169867, 25'd4260146, -25'd1689368, 25'd4774302, -25'd2350425}, '{-25'd8006137, -25'd6096416, -25'd5068105, -25'd7198178, -25'd6610572, -25'd3452187, -25'd1322114, -25'd220352, -25'd5655711}, '{-25'd6463670, -25'd4039794, -25'd7859235, -25'd2130073, -25'd3084933, -25'd8006137, -25'd7638883, -25'd1762819, 25'd146902}, '{-25'd7198178, 25'd0, -25'd1395565, -25'd6977825, -25'd3672540, -25'd4407048, -25'd2644229, -25'd1542467, -25'd6830924}}, '{'{25'd2717679, 25'd4113244, -25'd1248664, -25'd2423876, 25'd3672540, 25'd3378737, -25'd1395565, 25'd3231835, 25'd3452187}, '{-25'd734508, -25'd1322114, -25'd2497327, 25'd5068105, -25'd1101762, 25'd367254, 25'd2570778, 25'd293803, 25'd4847752}, '{-25'd293803, -25'd2570778, -25'd293803, 25'd2056622, 25'd3892892, 25'd440705, 25'd5215006, -25'd2423876, 25'd4260146}, '{-25'd3525638, 25'd1836270, 25'd3011483, 25'd1909721, 25'd2276975, 25'd2350425, 25'd146902, 25'd440705, 25'd3158384}, '{25'd3525638, 25'd2791130, -25'd2644229, 25'd2276975, 25'd4407048, -25'd1983171, 25'd5655711, 25'd6390219, 25'd4260146}, '{25'd5361908, 25'd3525638, 25'd2203524, -25'd1836270, 25'd514156, -25'd2864581, -25'd734508, 25'd3084933, 25'd4333597}, '{-25'd2276975, -25'd1395565, -25'd1248664, -25'd6830924, 25'd1542467, -25'd5729162, 25'd73451, -25'd1615917, -25'd8079587}, '{-25'd4627400, -25'd1689368, -25'd3892892, -25'd5068105, -25'd6830924, -25'd2350425, -25'd7124727, -25'd7712333, 25'd73451}, '{25'd1762819, -25'd440705, -25'd4553949, -25'd7345079, -25'd2938032, -25'd7418530, -25'd2791130, -25'd8006137, -25'd7565432}}},
    '{'{'{25'd3282472, 25'd3619135, -25'd2019983, -25'd1767485, 25'd336664, -25'd2314563, -25'd2146231, 25'd1893734, -25'd4587044}, '{25'd1178323, 25'd0, 25'd4713293, -25'd2062066, 25'd168332, -25'd715410, 25'd252498, -25'd4713293, -25'd3997882}, '{25'd4502878, 25'd1893734, -25'd1641236, -25'd294581, -25'd757493, 25'd2230397, 25'd2524978, 25'd1304572, 25'd420830}, '{25'd3577052, -25'd4124131, -25'd1346655, 25'd2440812, 25'd2693310, -25'd3619135, -25'd4797459, 25'd2861642, -25'd2693310}, '{25'd2062066, -25'd4292463, -25'd3450804, -25'd4208297, 25'd2945808, 25'd715410, 25'd3913716, 25'd3072057, -25'd336664}, '{25'd3324555, -25'd4755376, 25'd2819559, 25'd2146231, 25'd673328, 25'd2861642, -25'd841659, 25'd4208297, 25'd883742}, '{25'd2230397, -25'd1220406, 25'd3198306, 25'd4166214, -25'd3114140, -25'd3577052, -25'd3913716, 25'd336664, -25'd3324555}, '{25'd4502878, 25'd4713293, 25'd2861642, 25'd547079, 25'd3282472, 25'd0, -25'd4124131, 25'd1767485, -25'd1809568}, '{-25'd3240389, 25'd1220406, -25'd1262489, -25'd2777476, -25'd2482895, 25'd4166214, -25'd1977900, 25'd1809568, -25'd378747}}, '{'{-25'd2524978, -25'd378747, -25'd4587044, 25'd2651227, -25'd252498, 25'd3577052, 25'd84166, 25'd4208297, 25'd1009991}, '{-25'd4166214, -25'd1851651, -25'd84166, 25'd4166214, 25'd1388738, -25'd1767485, 25'd1178323, -25'd1725402, 25'd2146231}, '{-25'd1346655, 25'd2104149, 25'd3787467, -25'd2230397, 25'd3577052, -25'd3282472, 25'd3324555, -25'd2188314, -25'd2314563}, '{25'd3114140, -25'd4544961, -25'd883742, 25'd3156223, -25'd4502878, -25'd4713293, -25'd841659, -25'd2019983, -25'd2482895}, '{25'd3703301, 25'd1262489, -25'd631245, -25'd252498, 25'd715410, 25'd2819559, -25'd4334546, 25'd3997882, 25'd925825}, '{-25'd2019983, -25'd2482895, -25'd2987891, 25'd799576, 25'd420830, 25'd4166214, -25'd378747, -25'd3871633, -25'd547079}, '{-25'd4166214, -25'd2693310, 25'd2567061, -25'd1009991, -25'd2903725, 25'd504996, 25'd2272480, 25'd757493, 25'd2693310}, '{-25'd4376629, 25'd4502878, 25'd3787467, -25'd4208297, -25'd3408721, -25'd126249, 25'd1346655, -25'd1767485, 25'd1557070}, '{-25'd1052074, 25'd2861642, 25'd4418712, -25'd2019983, -25'd1557070, 25'd294581, 25'd504996, 25'd4587044, 25'd3114140}}, '{'{-25'd1683319, -25'd3240389, -25'd673328, 25'd2735393, -25'd4460795, -25'd3072057, -25'd1809568, -25'd3198306, 25'd3450804}, '{25'd925825, 25'd2567061, 25'd3534970, 25'd2356646, -25'd3198306, -25'd210415, 25'd4713293, 25'd3577052, 25'd2356646}, '{-25'd3661218, -25'd42083, -25'd3534970, 25'd3072057, 25'd1136240, 25'd4292463, -25'd2062066, -25'd1009991, 25'd3787467}, '{25'd84166, 25'd925825, 25'd3366638, -25'd1262489, 25'd1178323, 25'd1977900, -25'd42083, 25'd4039965, 25'd4502878}, '{-25'd4713293, -25'd3661218, -25'd1052074, 25'd3324555, 25'd5344537, 25'd1809568, 25'd4292463, 25'd4671210, 25'd4124131}, '{-25'd3029974, -25'd2019983, -25'd1557070, 25'd631245, -25'd799576, 25'd3955799, 25'd4376629, -25'd210415, 25'd883742}, '{-25'd925825, 25'd4124131, 25'd2735393, 25'd2272480, 25'd1557070, -25'd1052074, 25'd841659, -25'd1388738, -25'd2945808}, '{25'd3745384, 25'd2903725, 25'd2945808, 25'd4166214, 25'd4671210, 25'd2356646, -25'd1809568, -25'd4208297, -25'd1851651}, '{-25'd2314563, 25'd2524978, -25'd967908, 25'd1767485, -25'd3156223, 25'd2987891, -25'd2819559, -25'd799576, 25'd504996}}},
    '{'{'{-25'd2634970, 25'd4162489, 25'd4582557, -25'd916511, -25'd4620745, -25'd114564, 25'd649196, 25'd1527519, 25'd3742421}, '{25'd878323, 25'd2787722, -25'd2711346, 25'd3589669, -25'd2023962, 25'd1374767, -25'd458256, 25'd3666045, 25'd4315241}, '{25'd3971549, 25'd2176714, -25'd4200677, 25'd3131414, -25'd4391617, -25'd801947, 25'd229128, 25'd1222015, 25'd1489331}, '{-25'd1871211, -25'd954699, -25'd840135, -25'd2749534, -25'd2176714, -25'd3933361, -25'd3475105, -25'd2787722, -25'd2482218}, '{-25'd3245978, -25'd3093226, 25'd3016850, 25'd1680271, -25'd1794835, 25'd1412955, 25'd4773496, -25'd2711346, -25'd4811684}, '{-25'd4047925, 25'd4009737, -25'd954699, -25'd3475105, -25'd190940, -25'd4238865, 25'd2176714, 25'd916511, -25'd4849872}, '{25'd2023962, -25'd2749534, 25'd1489331, 25'd343692, -25'd152752, -25'd190940, -25'd3666045, -25'd1489331, 25'd992887}, '{25'd496444, -25'd2482218, 25'd1794835, 25'd3284166, -25'd3016850, 25'd1947587, -25'd2634970, 25'd878323, -25'd2940474}, '{-25'd2214902, -25'd4697121, 25'd2673158, 25'd2367654, -25'd2634970, -25'd4086113, -25'd4544369, -25'd4467993, -25'd2825910}}, '{'{-25'd4620745, -25'd840135, 25'd114564, -25'd3933361, -25'd114564, 25'd2138526, -25'd4811684, -25'd3780609, 25'd3895173}, '{-25'd2214902, -25'd572820, -25'd1183827, -25'd4506181, -25'd2864098, 25'd114564, -25'd3513293, 25'd1718459, -25'd3398729}, '{25'd114564, 25'd1336579, -25'd1909399, 25'd152752, -25'd725571, 25'd1489331, 25'd1833023, -25'd3436917, -25'd2100338}, '{-25'd458256, -25'd76376, 25'd2100338, -25'd1183827, 25'd3666045, 25'd725571, 25'd4009737, -25'd2444030, -25'd611008}, '{-25'd1489331, 25'd458256, -25'd2291278, -25'd2596782, 25'd2596782, 25'd267316, 25'd4506181, 25'd1947587, 25'd3895173}, '{-25'd2214902, 25'd3207790, 25'd2214902, -25'd916511, -25'd458256, -25'd3933361, 25'd4353429, 25'd2673158, -25'd114564}, '{-25'd3322354, 25'd4086113, 25'd4620745, -25'd152752, -25'd2444030, -25'd305504, 25'd4467993, 25'd190940, 25'd2558594}, '{-25'd3513293, 25'd4735308, -25'd3436917, -25'd4047925, -25'd4277053, -25'd38188, -25'd3513293, 25'd4544369, -25'd878323}, '{25'd2405842, -25'd3704233, 25'd4124301, -25'd3627857, 25'd3475105, -25'd2864098, -25'd3360542, 25'd4849872, 25'd2749534}}, '{'{-25'd2864098, -25'd1069263, -25'd4086113, 25'd2558594, 25'd1565707, -25'd1489331, -25'd1145639, 25'd4391617, -25'd649196}, '{25'd1909399, -25'd38188, -25'd3245978, -25'd2902286, -25'd2176714, 25'd611008, 25'd1107451, 25'd725571, 25'd1336579}, '{-25'd2902286, -25'd3513293, -25'd1145639, -25'd3627857, -25'd4124301, -25'd2176714, 25'd3169602, 25'd76376, 25'd3245978}, '{25'd611008, 25'd4047925, -25'd420068, -25'd114564, 25'd4277053, -25'd1069263, -25'd534632, -25'd2634970, -25'd2405842}, '{25'd3131414, 25'd3284166, 25'd3475105, 25'd3016850, -25'd2520406, 25'd1871211, -25'd4773496, -25'd3627857, 25'd4544369}, '{25'd1145639, -25'd3933361, 25'd38188, -25'd2673158, -25'd3780609, 25'd1603895, 25'd38188, 25'd1298391, 25'd3818797}, '{25'd1947587, 25'd458256, 25'd840135, 25'd1718459, -25'd992887, -25'd267316, 25'd2367654, -25'd1107451, 25'd1680271}, '{25'd3895173, -25'd2749534, 25'd420068, -25'd2787722, -25'd4506181, -25'd1222015, -25'd4047925, 25'd3818797, -25'd572820}, '{-25'd1565707, -25'd3207790, 25'd267316, 25'd4849872, -25'd2520406, 25'd3169602, 25'd1565707, 25'd1833023, -25'd3131414}}},
    '{'{'{-25'd1420911, 25'd2325127, -25'd3014054, -25'd1463969, -25'd4865544, 25'd1937606, 25'd1679259, -25'd4262733, 25'd3272401}, '{25'd2712648, 25'd2712648, -25'd4176617, 25'd2239011, 25'd3444633, 25'd215290, 25'd2798764, 25'd1808432, 25'd3487691}, '{-25'd5210007, -25'd2109838, -25'd1937606, 25'd1593143, 25'd1851490, -25'd5123891, -25'd3272401, -25'd2152896, 25'd3832154}, '{-25'd1463969, 25'd1894548, 25'd2970996, -25'd731984, 25'd1593143, 25'd602811, -25'd3100170, -25'd4521081, 25'd2712648}, '{-25'd2798764, -25'd516695, -25'd2884880, -25'd2195953, -25'd301405, -25'd4994718, -25'd5511413, -25'd4305791, -25'd5425297}, '{-25'd3487691, -25'd2152896, 25'd3918270, 25'd4564139, -25'd818100, -25'd2282069, 25'd2368185, -25'd2755706, -25'd1377853}, '{25'd3918270, -25'd4564139, 25'd5037776, 25'd4693312, -25'd861158, -25'd3918270, -25'd2841822, 25'd4176617, -25'd5468355}, '{25'd4908602, -25'd3789096, 25'd1593143, 25'd4133559, -25'd473637, 25'd1593143, 25'd818100, -25'd4004386, -25'd818100}, '{-25'd3444633, 25'd3401575, 25'd3746038, 25'd4865544, -25'd1593143, -25'd4779428, -25'd5511413, -25'd2325127, -25'd1033390}}, '{'{-25'd1076448, -25'd3487691, -25'd2841822, 25'd3315459, 25'd4693312, -25'd1550085, 25'd731984, 25'd775042, -25'd2411243}, '{-25'd5296123, -25'd43058, -25'd4521081, -25'd3014054, 25'd0, -25'd4478023, -25'd4650254, -25'd3616865, -25'd645869}, '{-25'd3229343, -25'd2841822, -25'd5425297, 25'd3358517, -25'd1420911, 25'd2927938, 25'd4176617, -25'd4348849, 25'd1593143}, '{-25'd3573807, -25'd4693312, 25'd86116, -25'd3315459, 25'd2755706, -25'd2669590, -25'd4004386, 25'd1377853, 25'd861158}, '{-25'd1076448, -25'd2626533, 25'd2497359, 25'd4478023, 25'd4693312, -25'd559753, -25'd5511413, 25'd1291737, -25'd1593143}, '{-25'd1679259, 25'd1420911, -25'd2454301, 25'd5382239, -25'd3186285, 25'd430579, -25'd1894548, 25'd4736370, 25'd2066780}, '{-25'd1550085, 25'd3702980, 25'd2454301, -25'd1420911, 25'd5339181, 25'd4391907, -25'd1679259, 25'd301405, -25'd1291737}, '{25'd3143227, 25'd1765374, 25'd4779428, -25'd2282069, 25'd2927938, -25'd215290, 25'd2282069, -25'd1291737, -25'd4564139}, '{25'd1550085, 25'd4779428, -25'd3229343, -25'd3014054, -25'd387521, 25'd3057112, 25'd2368185, -25'd1076448, 25'd2798764}}, '{'{25'd2023722, -25'd1593143, -25'd1377853, -25'd2884880, 25'd775042, 25'd3444633, 25'd4219675, 25'd2282069, -25'd258347}, '{25'd1722316, -25'd2497359, -25'd129174, -25'd3057112, 25'd430579, -25'd1420911, 25'd775042, 25'd3530749, -25'd645869}, '{25'd1119506, -25'd5425297, -25'd947274, -25'd1894548, 25'd1291737, -25'd1851490, -25'd3315459, -25'd1507027, -25'd43058}, '{-25'd3186285, -25'd43058, 25'd516695, -25'd4951660, 25'd2970996, -25'd3143227, -25'd3530749, 25'd2755706, 25'd559753}, '{-25'd861158, -25'd947274, 25'd3143227, -25'd1593143, 25'd3487691, 25'd904216, 25'd2066780, -25'd2755706, -25'd2712648}, '{25'd5166949, -25'd1248679, 25'd4004386, -25'd86116, -25'd3875212, -25'd129174, 25'd688927, 25'd4391907, -25'd5037776}, '{25'd1463969, -25'd947274, -25'd2884880, 25'd1980664, -25'd2195953, -25'd4951660, -25'd1420911, 25'd3358517, 25'd2368185}, '{25'd5080833, -25'd4047444, 25'd301405, 25'd4736370, -25'd2583475, -25'd4478023, -25'd5511413, -25'd3702980, 25'd1722316}, '{-25'd2454301, 25'd1550085, 25'd2970996, 25'd1119506, -25'd1463969, 25'd4348849, -25'd4176617, 25'd4521081, -25'd775042}}},
    '{'{'{25'd3585482, 25'd4860319, 25'd2669192, 25'd119516, -25'd876451, 25'd756935, -25'd4501771, 25'd3784675, -25'd2908224}, '{25'd438226, -25'd1115483, -25'd3426127, 25'd4541610, 25'd3744836, 25'd3346449, 25'd995967, 25'd2031773, -25'd2669192}, '{-25'd796774, 25'd2948063, -25'd4461933, 25'd318709, -25'd677258, -25'd3585482, 25'd239032, 25'd4700965, 25'd1314677}, '{25'd1354515, -25'd1752902, -25'd3983868, -25'd239032, -25'd1115483, -25'd4939997, 25'd717096, 25'd3505804, -25'd3824514}, '{-25'd278871, 25'd39839, 25'd2748869, -25'd239032, -25'd637419, -25'd2310644, 25'd597580, -25'd358548, 25'd119516}, '{25'd1713063, -25'd3067579, 25'd478064, 25'd3306611, 25'd1155322, -25'd2748869, 25'd39839, 25'd4581449, -25'd3744836}, '{-25'd4382255, 25'd5059513, -25'd1513870, 25'd4382255, -25'd4621287, 25'd2589514, -25'd4143223, 25'd5019674, -25'd1234999}, '{25'd3306611, -25'd677258, -25'd717096, -25'd2908224, -25'd3585482, -25'd2788708, -25'd3306611, -25'd3226933, 25'd2071612}, '{25'd4422094, 25'd3027740, -25'd1952096, 25'd2589514, -25'd2151289, 25'd3704998, -25'd1991934, -25'd199193, 25'd4661126}}, '{'{-25'd557742, -25'd4342417, 25'd2469998, 25'd995967, 25'd2151289, 25'd358548, 25'd3744836, 25'd3147256, -25'd2589514}, '{-25'd79677, -25'd1832579, -25'd318709, -25'd159355, -25'd4143223, -25'd159355, -25'd2828547, 25'd3904191, -25'd3625320}, '{25'd4501771, -25'd1832579, -25'd2071612, -25'd1274838, -25'd876451, -25'd1354515, 25'd4979835, -25'd318709, 25'd2589514}, '{-25'd916290, -25'd239032, -25'd3744836, -25'd1155322, 25'd0, -25'd2191128, 25'd3864352, -25'd39839, 25'd2908224}, '{25'd2350482, -25'd4222900, -25'd119516, 25'd3505804, -25'd756935, 25'd3465966, 25'd4541610, 25'd3904191, 25'd3067579}, '{25'd4222900, 25'd4661126, -25'd517903, 25'd4222900, 25'd3704998, 25'd557742, 25'd2191128, 25'd2629353, 25'd2111450}, '{-25'd3465966, 25'd5059513, 25'd995967, 25'd717096, -25'd3147256, -25'd1832579, 25'd1752902, -25'd2709031, 25'd119516}, '{-25'd3187095, -25'd4422094, 25'd3067579, 25'd438226, -25'd677258, -25'd4621287, 25'd2111450, -25'd1274838, 25'd2071612}, '{-25'd2350482, -25'd3067579, -25'd1832579, -25'd3266772, 25'd3226933, 25'd0, -25'd278871, -25'd4541610, 25'd2709031}}, '{'{25'd1035806, -25'd4262739, -25'd2788708, -25'd1713063, 25'd3944030, -25'd1394354, -25'd2629353, -25'd637419, 25'd1075644}, '{25'd3904191, -25'd398387, 25'd3545643, -25'd2111450, 25'd3665159, -25'd517903, 25'd2230966, 25'd2868385, -25'd4023707}, '{-25'd3027740, 25'd1593547, 25'd4103384, 25'd4740803, 25'd1314677, 25'd119516, 25'd478064, 25'd3465966, 25'd79677}, '{25'd478064, 25'd4063546, -25'd2828547, 25'd4143223, 25'd2669192, -25'd119516, -25'd517903, -25'd3545643, 25'd1314677}, '{-25'd1035806, 25'd836612, -25'd3187095, 25'd2509837, 25'd1314677, 25'd3585482, 25'd4700965, 25'd2111450, 25'd2868385}, '{-25'd1593547, 25'd1593547, 25'd3824514, 25'd1752902, -25'd3904191, 25'd1633386, -25'd3147256, 25'd4621287, 25'd4183062}, '{25'd1314677, -25'd2191128, -25'd4541610, 25'd3625320, 25'd3465966, 25'd3226933, -25'd4143223, -25'd79677, -25'd2111450}, '{-25'd1832579, -25'd3505804, -25'd3386288, 25'd2908224, -25'd318709, 25'd4621287, -25'd3744836, -25'd2908224, 25'd1394354}, '{25'd4860319, -25'd1792741, -25'd2509837, 25'd3306611, 25'd3625320, -25'd1713063, -25'd2868385, -25'd2589514, -25'd1633386}}},
    '{'{'{-25'd1748028, 25'd635647, 25'd516463, -25'd3416601, -25'd1469933, -25'd1152110, 25'd2145307, -25'd2741226, 25'd2224763}, '{25'd2979594, 25'd953470, -25'd1986396, 25'd2542587, -25'd834286, -25'd2820682, -25'd158912, -25'd3297417, 25'd2145307}, '{-25'd2463131, 25'd2860410, 25'd2542587, -25'd3575512, 25'd3456329, 25'd1152110, 25'd357551, 25'd3575512, 25'd476735}, '{-25'd2542587, 25'd1112382, -25'd993198, 25'd4370071, 25'd2185035, -25'd2423403, -25'd2900138, 25'd715102, -25'd4290615}, '{-25'd2065852, -25'd1469933, -25'd3178233, 25'd913742, -25'd3535784, 25'd4449527, 25'd1271293, -25'd3178233, -25'd5085173}, '{-25'd2820682, -25'd2780954, 25'd3813880, -25'd3734424, -25'd2979594, 25'd4131703, 25'd2582315, -25'd4846806, -25'd4330343}, '{-25'd4886534, 25'd2820682, -25'd4886534, 25'd993198, 25'd357551, -25'd2502859, -25'd1946668, -25'd4727622, 25'd2026124}, '{25'd1787756, -25'd4091975, 25'd1231565, 25'd1708300, 25'd2185035, 25'd2105580, 25'd158912, 25'd4211159, 25'd2502859}, '{25'd3734424, -25'd4648166, 25'd2860410, 25'd3734424, 25'd1549389, 25'd2979594, 25'd3893336, -25'd4608438, 25'd476735}}, '{'{25'd1509661, -25'd4886534, 25'd238367, -25'd1271293, -25'd4727622, 25'd595919, -25'd1430205, -25'd953470, 25'd437007}, '{25'd1906940, 25'd4012519, 25'd4052247, -25'd317823, 25'd2820682, -25'd635647, -25'd1906940, -25'd3257689, -25'd1549389}, '{25'd2463131, -25'd1906940, -25'd1946668, 25'd4012519, -25'd79456, -25'd754830, -25'd794558, -25'd2741226, -25'd3654968}, '{-25'd4370071, -25'd913742, -25'd5005717, 25'd3257689, 25'd2582315, 25'd2542587, -25'd754830, 25'd4250887, -25'd675375}, '{25'd3337145, 25'd4489254, 25'd1311021, 25'd1589117, -25'd317823, -25'd1589117, -25'd2701498, -25'd4330343, -25'd4807078}, '{-25'd3933064, 25'd158912, 25'd913742, 25'd3654968, 25'd4687894, 25'd357551, -25'd3535784, -25'd2820682, 25'd2065852}, '{-25'd3416601, -25'd2741226, -25'd4449527, 25'd1469933, -25'd3893336, 25'd913742, -25'd2145307, 25'd1231565, 25'd1906940}, '{-25'd1271293, -25'd1668572, -25'd3098777, -25'd2383675, 25'd1032926, 25'd1628845, 25'd3178233, -25'd516463, -25'd3813880}, '{25'd3496057, -25'd79456, 25'd2979594, -25'd2979594, -25'd3774152, -25'd437007, -25'd1350749, -25'd1628845, -25'd4250887}}, '{'{-25'd3933064, 25'd4727622, -25'd4449527, -25'd3416601, 25'd1906940, 25'd3774152, 25'd2304219, 25'd3535784, -25'd1032926}, '{-25'd2105580, -25'd4965989, 25'd119184, 25'd1827484, 25'd1549389, 25'd2622042, 25'd278095, -25'd119184, -25'd3217961}, '{25'd2264491, -25'd3217961, -25'd4290615, -25'd834286, -25'd4489254, 25'd4171431, -25'd4648166, -25'd1628845, 25'd1708300}, '{-25'd1827484, -25'd2582315, 25'd2979594, -25'd3456329, -25'd3376873, -25'd4211159, 25'd4608438, 25'd993198, -25'd675375}, '{25'd3496057, 25'd3575512, 25'd913742, 25'd4250887, -25'd238367, 25'd2622042, -25'd2780954, -25'd4211159, 25'd357551}, '{-25'd794558, -25'd3774152, -25'd4727622, 25'd1549389, 25'd238367, 25'd3575512, -25'd1748028, 25'd1390477, 25'd4409799}, '{-25'd1430205, -25'd4528982, -25'd2741226, 25'd3019322, 25'd2741226, -25'd1628845, 25'd4171431, -25'd158912, 25'd1549389}, '{-25'd1986396, 25'd1469933, -25'd2026124, -25'd238367, -25'd1708300, -25'd4409799, -25'd2780954, -25'd3217961, 25'd3138505}, '{-25'd3972792, -25'd238367, 25'd1152110, 25'd1946668, 25'd2145307, 25'd2502859, -25'd1787756, -25'd675375, 25'd4608438}}}
};
