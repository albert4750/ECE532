localparam bit signed [0:26][19:0] Output4 = '{20'd106, -20'd8, 20'd199, -20'd217, 20'd90, -20'd237, 20'd12, -20'd127, 20'd138, -20'd29, -20'd65, 20'd50, -20'd142, -20'd8, -20'd133, -20'd229, 20'd121, -20'd232, -20'd81, 20'd2, 20'd258, 20'd51, -20'd36, -20'd155, -20'd134, -20'd17, -20'd111};
