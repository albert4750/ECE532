localparam bit signed [0:146][7:0] Input8 = '{9, 46, 60, -52, 101, 29, -19, -53, 108, 105, -15, 24, -69, 72, 15, 54, 32, 108, 126, 80, 114, -13, -20, -14, -15, -117, -113, -103, -107, 22, 81, 92, 122, -37, -20, 72, -37, 92, 103, -21, -25, -29, 30, 116, 41, 118, 9, -10, -76, -85, -47, 50, 16, -64, -102, 7, 54, -46, 58, -53, -71, 58, 76, -115, 72, 104, -110, 17, 42, -84, 98, 75, -41, -58, 78, -82, -74, 50, -85, -63, 78, -27, -122, -7, 47, 44, -119, -125, 9, -5, 116, 123, -94, 94, -127, -90, 78, 80, -34, 50, 13, -42, -82, 99, -41, -91, -35, 109, 106, -38, -46, 86, -122, -54, 43, -127, 73, 90, 48, -49, 17, -109, 126, 19, -63, 27, 115, 100, 35, -119, 105, -115, 53, -58, 88, -118, -7, -85, -27, 5, 40, 116, -113, -114, 85, -128, -93};
