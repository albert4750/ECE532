localparam bit signed [0:2][0:26][19:0] Input8 = '{
    '{20'd73, 20'd53, 20'd69, 20'd33, 20'd7, -20'd3, -20'd34, -20'd56, 20'd118, -20'd44, 20'd7, 20'd67, 20'd85, 20'd91, -20'd20, -20'd61, -20'd26, -20'd44, -20'd57, -20'd45, 20'd95, -20'd128, 20'd5, -20'd37, -20'd21, 20'd30, 20'd73},
    '{20'd83, -20'd121, 20'd21, 20'd101, 20'd92, 20'd8, 20'd43, -20'd82, -20'd128, -20'd24, 20'd51, -20'd90, -20'd39, -20'd54, 20'd115, 20'd98, -20'd5, -20'd41, -20'd32, -20'd45, -20'd102, 20'd78, -20'd96, -20'd13, 20'd70, -20'd31, 20'd44},
    '{-20'd69, -20'd71, 20'd50, 20'd45, 20'd105, 20'd4, 20'd57, -20'd35, -20'd37, 20'd17, 20'd35, 20'd66, 20'd20, 20'd45, 20'd57, 20'd79, -20'd9, 20'd36, -20'd23, 20'd62, -20'd124, 20'd113, 20'd114, 20'd77, 20'd30, -20'd19, -20'd41}
};
