logic signed [7:0] convolve19_weight[4][8][3][3] = '{
    '{
        '{'{120, 31, -42}, '{-71, 114, -105}, '{-4, -60, -64}},
        '{'{17, 70, -60}, '{75, 96, 80}, '{2, 122, 74}},
        '{'{39, 126, 38}, '{54, 124, -25}, '{125, 119, 0}},
        '{'{-119, -53, 44}, '{-76, 81, -28}, '{-23, 47, 69}},
        '{'{105, -80, 38}, '{-92, 4, 123}, '{113, 75, -89}},
        '{'{93, 107, 62}, '{45, 75, -86}, '{32, 1, 108}},
        '{'{47, 34, -86}, '{-86, -20, 74}, '{42, 124, 104}},
        '{'{-82, 103, 79}, '{-19, 90, -23}, '{-88, -20, -16}}
    },
    '{
        '{'{-48, 43, -36}, '{64, -65, -84}, '{-3, 2, -106}},
        '{'{-4, 24, 44}, '{-45, 94, 77}, '{7, 83, 99}},
        '{'{-75, 117, -66}, '{29, 84, -120}, '{74, -87, 34}},
        '{'{46, 61, 75}, '{125, 72, -11}, '{-73, 85, 116}},
        '{'{-60, -81, -121}, '{120, -72, -43}, '{-42, -58, -109}},
        '{'{43, -58, -32}, '{123, -27, -42}, '{-23, -107, 116}},
        '{'{11, 43, -61}, '{96, 29, 21}, '{81, -59, 111}},
        '{'{91, -127, 33}, '{40, -21, -25}, '{121, 43, -77}}
    },
    '{
        '{'{101, -34, 82}, '{54, 79, 124}, '{-77, 45, 104}},
        '{'{-35, 4, 56}, '{48, -8, 106}, '{20, -112, -75}},
        '{'{85, 66, 20}, '{109, 56, 24}, '{-85, -44, 109}},
        '{'{63, -113, -31}, '{-104, -40, -24}, '{-37, -67, 3}},
        '{'{19, 12, -14}, '{-84, -54, 9}, '{63, 92, -11}},
        '{'{46, 95, 87}, '{13, -59, 45}, '{104, 7, -87}},
        '{'{-18, 16, 50}, '{-89, -93, -22}, '{-100, -11, -47}},
        '{'{-91, -127, 81}, '{-98, -94, -12}, '{-125, 33, 43}}
    },
    '{
        '{'{-39, -127, -30}, '{56, -79, -25}, '{-88, -46, -87}},
        '{'{-74, 85, 47}, '{-36, -1, 65}, '{-87, -90, 12}},
        '{'{79, 28, -103}, '{123, 114, -75}, '{86, 63, -37}},
        '{'{-51, 33, 78}, '{-11, 8, 68}, '{-82, -10, -43}},
        '{'{45, 92, -106}, '{-114, -128, 50}, '{101, 54, 50}},
        '{'{9, -95, 116}, '{-88, 40, 115}, '{7, 26, 29}},
        '{'{50, 57, -111}, '{-2, -118, -85}, '{62, 97, 65}},
        '{'{102, -3, -109}, '{93, 6, -123}, '{68, 66, 119}}
    }
};
