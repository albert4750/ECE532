logic signed [7:0] convolve7_weight[4][8][3][3] = '{
    '{
        '{'{71, -68, -104}, '{32, -20, -89}, '{-12, -24, -2}},
        '{'{-17, -12, 100}, '{106, -112, 52}, '{90, 104, 80}},
        '{'{-82, 96, -34}, '{-44, -105, 15}, '{44, -45, -9}},
        '{'{-73, -30, 27}, '{-83, 98, -47}, '{87, 27, -51}},
        '{'{48, 87, -34}, '{5, -7, 103}, '{97, -15, 98}},
        '{'{-100, 116, -63}, '{-60, 85, 72}, '{124, -14, 33}},
        '{'{-10, 99, -80}, '{-29, 89, -59}, '{65, -29, -57}},
        '{'{-127, 1, 71}, '{25, -28, -51}, '{-20, 50, 27}}
    },
    '{
        '{'{-32, -85, -109}, '{-30, -83, -28}, '{-48, -16, 106}},
        '{'{-7, 43, 67}, '{-120, 83, 46}, '{-64, -12, 20}},
        '{'{-32, 98, -21}, '{5, -43, -104}, '{-126, 125, 125}},
        '{'{71, -20, 75}, '{115, -100, -10}, '{-33, -63, 80}},
        '{'{-14, 82, 14}, '{-107, -17, -17}, '{69, -95, -22}},
        '{'{2, -101, 104}, '{-9, 19, 15}, '{-57, 108, -99}},
        '{'{35, 97, -80}, '{49, -48, 56}, '{-65, 88, 58}},
        '{'{5, -77, 122}, '{-67, -22, 83}, '{-111, -83, 96}}
    },
    '{
        '{'{-66, -106, 97}, '{-26, 9, -123}, '{-52, -67, 42}},
        '{'{119, 16, -69}, '{-111, 68, -68}, '{25, 14, -19}},
        '{'{-67, 53, -47}, '{-99, 70, -100}, '{74, 5, 100}},
        '{'{100, -44, 55}, '{114, 50, -42}, '{53, -118, -85}},
        '{'{59, 30, -69}, '{14, 115, 48}, '{-8, -3, -72}},
        '{'{65, -24, 7}, '{69, 15, -9}, '{105, -76, -96}},
        '{'{-41, 78, 34}, '{-99, -77, 89}, '{53, -124, 64}},
        '{'{-5, 26, 84}, '{5, -6, -40}, '{-111, 68, -72}}
    },
    '{
        '{'{32, 113, -47}, '{-56, -55, 100}, '{31, -34, -55}},
        '{'{-20, 48, 99}, '{32, -114, -67}, '{-41, 32, -72}},
        '{'{28, 43, -31}, '{50, -82, -20}, '{-56, 37, -8}},
        '{'{-126, -111, 15}, '{67, -43, 112}, '{114, -35, -27}},
        '{'{-8, 22, 82}, '{-121, -73, 49}, '{-102, 120, 4}},
        '{'{-19, -39, -102}, '{60, 115, -17}, '{-45, -50, 18}},
        '{'{-7, -32, -37}, '{-92, -26, 20}, '{-1, 108, 3}},
        '{'{18, 77, -77}, '{-79, -97, 97}, '{18, -116, -17}}
    }
};
