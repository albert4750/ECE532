logic signed [7:0] convolve20_weight[4][8][3][3] = '{
    '{
        '{'{40, 104, 80}, '{-57, 40, -104}, '{87, 52, -6}},
        '{'{22, -87, -122}, '{-8, 78, -77}, '{39, 127, -104}},
        '{'{-97, 20, 18}, '{-93, 96, 84}, '{-40, 96, -37}},
        '{'{-84, 122, -28}, '{82, 22, 98}, '{31, 50, -110}},
        '{'{124, -50, -121}, '{-117, 63, 74}, '{57, -70, -90}},
        '{'{41, 86, 64}, '{-94, 81, 42}, '{52, -58, 3}},
        '{'{40, -5, -37}, '{76, 39, 85}, '{-103, -128, -21}},
        '{'{34, -3, 65}, '{-16, -85, 37}, '{110, -21, 89}}
    },
    '{
        '{'{87, -86, 115}, '{68, 52, 71}, '{-35, -127, -105}},
        '{'{87, -40, -39}, '{-59, 22, 113}, '{-48, -33, 112}},
        '{'{64, 114, 67}, '{-31, -97, 70}, '{-76, -64, -120}},
        '{'{-104, -58, -53}, '{68, -66, 117}, '{-27, -57, 119}},
        '{'{-103, 51, -86}, '{5, 37, 4}, '{124, 127, 62}},
        '{'{-86, 121, -116}, '{-112, 57, -59}, '{-115, -117, 86}},
        '{'{-22, -89, -128}, '{24, -16, 27}, '{-9, 30, 88}},
        '{'{92, 24, 127}, '{-2, -34, -7}, '{52, -18, 32}}
    },
    '{
        '{'{62, -67, 110}, '{99, -42, -81}, '{8, -125, -28}},
        '{'{52, 78, -68}, '{100, -69, 81}, '{59, 83, -40}},
        '{'{-40, -29, 114}, '{-63, 76, -44}, '{-121, -42, -84}},
        '{'{120, 79, -96}, '{-95, -51, 1}, '{-125, 39, 120}},
        '{'{62, -66, -28}, '{102, -101, 58}, '{-30, -19, 102}},
        '{'{47, 25, -48}, '{112, -14, 127}, '{73, 25, 64}},
        '{'{-113, 117, -48}, '{106, 125, -28}, '{-121, 23, 113}},
        '{'{-88, -90, -19}, '{-91, -15, -27}, '{68, 98, -42}}
    },
    '{
        '{'{60, 122, -79}, '{-98, 123, 97}, '{91, -57, 77}},
        '{'{89, 37, 31}, '{100, 122, 49}, '{47, -75, -25}},
        '{'{8, -110, 84}, '{-103, 39, 93}, '{-126, 104, 50}},
        '{'{81, -24, -25}, '{-31, -125, -102}, '{53, -17, 88}},
        '{'{63, 127, 127}, '{-15, 94, -13}, '{57, -63, -22}},
        '{'{-46, -57, 43}, '{-59, -70, 40}, '{-27, 19, -94}},
        '{'{85, 100, -40}, '{-34, 65, 0}, '{88, -19, -81}},
        '{'{-8, -124, -64}, '{36, -68, 50}, '{55, 84, -60}}
    }
};
