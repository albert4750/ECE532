localparam bit signed [0:46][15:0] Input9 = '{-16'd428, -16'd9750, 16'd11585, 16'd6007, -16'd29164, -16'd29488, -16'd27606, 16'd5618, 16'd16412, 16'd1434, 16'd2903, 16'd3252, -16'd26320, 16'd14274, -16'd6554, -16'd7415, -16'd25342, -16'd21132, 16'd31596, -16'd2327, 16'd13145, 16'd13692, -16'd7307, -16'd32156, -16'd28582, -16'd7100, 16'd25193, 16'd9738, -16'd12276, 16'd22120, 16'd10465, -16'd5723, -16'd12121, -16'd23648, 16'd25978, 16'd11553, -16'd23654, -16'd32669, 16'd23769, -16'd30414, 16'd26968, 16'd31954, 16'd22292, 16'd13022, 16'd32412, -16'd31160, 16'd21778};
