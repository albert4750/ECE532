localparam bit signed [0:46][15:0] Input6 = '{16'd31915, 16'd18131, 16'd11096, 16'd32326, -16'd24940, -16'd7290, 16'd3868, -16'd11661, 16'd4998, -16'd27838, 16'd16988, 16'd24540, 16'd3686, -16'd7323, -16'd12933, -16'd12603, -16'd19347, 16'd9545, -16'd32668, 16'd21174, -16'd23731, -16'd26731, 16'd22011, -16'd7521, 16'd20049, 16'd19491, -16'd7955, 16'd15603, 16'd14586, -16'd1656, 16'd23294, 16'd9497, -16'd16363, -16'd9811, 16'd17637, 16'd6102, -16'd7792, -16'd2919, 16'd25582, -16'd29577, 16'd9893, 16'd8063, 16'd30081, 16'd30085, 16'd18118, 16'd6540, -16'd29350};
