localparam bit signed [0:10][15:0] Output5 = '{16'd2781, -16'd19400, 16'd6759, 16'd7658, -16'd9018, 16'd735, -16'd17363, 16'd9366, 16'd4769, -16'd26849, 16'd18818};
