logic signed [7:0] convolve14_weight[4][8][3][3] = '{
    '{
        '{'{-115, 8, 6}, '{27, 37, 35}, '{-88, 26, -34}},
        '{'{76, 57, -83}, '{-48, -70, 23}, '{126, 114, 106}},
        '{'{72, 119, 118}, '{80, 117, -3}, '{-110, 74, 15}},
        '{'{102, -3, -40}, '{100, 111, -64}, '{3, 90, 20}},
        '{'{111, 47, 62}, '{-31, -104, 82}, '{-88, 9, -56}},
        '{'{71, 92, 111}, '{-87, -109, 86}, '{-61, 119, 78}},
        '{'{-1, -9, -62}, '{87, 107, -104}, '{-44, 35, -6}},
        '{'{46, -96, -94}, '{-86, -36, -91}, '{100, -46, -73}}
    },
    '{
        '{'{-22, -93, 103}, '{-29, -63, -35}, '{20, 101, -29}},
        '{'{-82, -30, -37}, '{-66, -66, 113}, '{123, -50, -22}},
        '{'{30, -37, -77}, '{-124, 68, 6}, '{105, -87, -125}},
        '{'{39, 108, -28}, '{27, 13, -84}, '{-128, -54, 93}},
        '{'{-50, 0, -128}, '{-32, -12, -117}, '{-99, 5, -59}},
        '{'{57, -98, -110}, '{-22, -112, -9}, '{-47, 75, -119}},
        '{'{9, 90, -52}, '{64, 103, 28}, '{118, -51, -41}},
        '{'{58, -7, 48}, '{27, -21, 25}, '{84, -17, -52}}
    },
    '{
        '{'{-104, -123, -94}, '{-52, 59, -85}, '{79, -69, -107}},
        '{'{100, 113, 126}, '{-20, -116, -16}, '{-30, 5, -108}},
        '{'{-4, 31, -30}, '{-105, -109, -43}, '{-81, 122, -122}},
        '{'{-60, 73, -104}, '{47, 32, 74}, '{90, 91, -112}},
        '{'{98, 22, -3}, '{-100, -100, -15}, '{78, -27, -39}},
        '{'{5, -62, 35}, '{75, 51, -51}, '{99, 56, 95}},
        '{'{94, -123, -99}, '{-37, 121, 53}, '{65, -67, 104}},
        '{'{26, -100, 103}, '{39, -31, -23}, '{47, -19, 32}}
    },
    '{
        '{'{-7, -124, 54}, '{0, -117, 51}, '{-29, 68, -102}},
        '{'{-113, 113, 92}, '{-22, 16, -12}, '{-58, 120, -33}},
        '{'{-126, 124, -111}, '{114, -63, 32}, '{97, 38, -60}},
        '{'{-34, -124, 123}, '{-49, -1, -107}, '{-7, -13, -26}},
        '{'{-118, -112, -126}, '{-82, 61, 46}, '{-18, -96, 103}},
        '{'{23, 61, 1}, '{-92, -39, -120}, '{-81, -37, -128}},
        '{'{35, -102, 62}, '{-17, 52, 106}, '{22, 31, 1}},
        '{'{-35, -125, -125}, '{-30, -12, 36}, '{42, -18, -108}}
    }
};
