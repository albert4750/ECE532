logic signed [15:0] layer1_weight[16][3][7][7] = '{
    '{
        '{'{-30036, 10799, 9845, 19648, 13123, -11525, -2365}, '{-665, 9225, 24275, -12011, 22258, 14116, -17833}, '{-17338, 15832, 6744, 19852, -18118, -15679, -538}, '{-13785, 10327, 18606, -8616, 2897, 26277, -15847}, '{-5299, 6216, -25847, 6036, -30605, -27696, 4851}, '{-24891, -14338, -30897, -25169, -30272, 15186, -8093}, '{10200, -847, 755, -31971, 17043, -29549, -17522}},
        '{'{-7769, 23840, -16447, 19721, -13639, 21119, 8736}, '{23071, 17098, -14092, 24727, 27299, -1538, -21045}, '{11122, -15177, 22556, 25378, 10368, -6016, 26532}, '{-9163, -26747, -12762, -29208, -7436, 28945, -1713}, '{12676, 18025, 27690, 13754, 14879, -11400, -12031}, '{30017, -4121, 28585, -6087, -18141, -20634, 27767}, '{15115, 8622, 23634, -12197, 30592, 27022, 19043}},
        '{'{-22987, -13428, -5511, -16470, -20396, 18635, -28348}, '{13062, 7108, -15313, 29311, -18444, 5251, 29644}, '{-25756, -23372, 14312, -28850, -23409, 18068, 11491}, '{-9286, -17641, 10959, 2957, 4469, -18603, -24016}, '{30001, 9797, -18263, -26973, 17856, -9121, 7365}, '{-4514, 8448, 22385, 3762, 29988, 26530, -7376}, '{-16547, -13949, 1634, 15914, -31795, -11920, -22553}}
    },
    '{
        '{'{-21611, -7991, 27007, -18944, 30602, -30350, -19925}, '{-19526, 3455, 22551, 22203, 28802, -26247, -10142}, '{24126, -23645, -1314, 30843, 10179, 23122, -18514}, '{19171, -9068, 4305, 18994, 5531, -9458, -983}, '{31802, -17727, 23588, -9462, 4182, 15403, -19608}, '{-6133, 15106, 307, -19376, -18400, -27466, 1152}, '{-9434, 8467, 5294, 13866, 13683, 17592, 2492}},
        '{'{-5656, 15949, 14622, -19176, -7555, 770, -16893}, '{-24482, 11490, 5995, 32013, 30576, -14040, -19128}, '{-29677, 12895, -28856, 17818, -26174, -11016, 24756}, '{26947, -9236, -24771, 20238, 8032, -17148, 8131}, '{-27923, -6005, 21500, 10838, -29235, -29831, -6547}, '{4939, 31416, 9744, -13160, -27747, -5995, 1134}, '{16409, 9680, -15428, -30855, 19318, -19339, 26045}},
        '{'{-18861, 2721, -22680, 17312, -17180, 5627, 27387}, '{22649, 5446, -32299, 10527, -24051, 18247, 1720}, '{5272, -15793, 6185, 18706, -16856, -4682, -16177}, '{-17653, 20646, -18321, 19805, -4103, 21633, 31455}, '{10102, -21716, 24792, -17027, 24600, -4029, 11218}, '{-27665, 24323, 2282, -31028, 22502, -20189, -26922}, '{13310, 15037, -12603, -29993, -13781, -2016, -9205}}
    },
    '{
        '{'{-18840, -26412, 1162, 14006, -4117, 30117, -16771}, '{32412, 623, -536, -23806, 30235, -12333, 1241}, '{10903, 25397, -28365, -15186, -2924, -13387, 5661}, '{-16829, -21981, -15577, 28041, -30647, 12585, 31639}, '{-8317, -28882, 8922, -10318, -17556, -22781, 18207}, '{15113, 28042, 28187, 12717, -16185, 1447, -27587}, '{10581, 29537, 27692, -21726, 10146, -27560, -26591}},
        '{'{14981, 30952, -27905, 22564, 18176, 17867, 14626}, '{-24379, -31874, 30645, 21758, 15440, -2626, 136}, '{-5955, 6273, 26833, -6800, 14627, -19080, -29349}, '{-16216, -26764, 2852, 12464, 9753, -11965, 24423}, '{25084, -17629, 3186, -10466, -11235, -14607, 19745}, '{8338, 21777, 20701, -18092, -11779, -30206, -10171}, '{30053, -7284, 4652, -19595, -5379, 13634, -4497}},
        '{'{22619, -21163, 423, 28199, 32715, -4458, 28062}, '{28305, 23238, 967, 4370, 9052, -10197, 21587}, '{433, -19671, -10147, 29870, -14955, 28873, 12121}, '{-13838, -1568, -18469, -16055, -12772, -16405, -7983}, '{23145, 30650, 3968, -8234, -449, -31728, -26518}, '{24740, -7586, -25064, -25996, 5311, 9411, -6861}, '{12424, -23624, 29531, -5027, 6011, 19182, 29783}}
    },
    '{
        '{'{8352, -30573, -28088, 22983, -7081, 19469, -710}, '{22097, 5240, -22668, 27575, -17600, 10955, 732}, '{21412, 24857, 13088, -8790, -20722, -11818, -23268}, '{7444, -46, 19780, 13846, 21731, -9350, 16979}, '{647, -20536, -15811, 6797, 5637, 24832, -4984}, '{11471, 14799, -75, 5259, 9220, 6567, 4444}, '{19373, 29978, 586, -18636, 21486, -25167, -4901}},
        '{'{-21709, -32029, -3223, -11502, -4747, -27358, 15923}, '{16030, -15947, -28870, -4181, -14537, -23044, 17404}, '{-9454, -31827, -5289, -7743, -21178, 21994, -21451}, '{-23760, -930, -14277, -18096, -6502, -2436, -12125}, '{-20934, -15439, 29802, -24375, 23852, -14579, 15225}, '{-30906, 8742, 3751, 9864, 31757, 18424, -31865}, '{-2352, -17416, 31254, -7688, -8369, -18471, -26872}},
        '{'{-20765, -24826, -9007, 9671, 31188, 5593, -16446}, '{-2500, 29072, 19512, 7026, 3821, -13673, -24296}, '{-31740, 2660, 29676, -30415, -5801, -10722, -25034}, '{-8039, -4332, -8863, -5787, -21831, 12695, -613}, '{-31715, -13407, -10893, 3893, -30089, -21581, -27818}, '{-1546, 28679, -30103, -13327, -1911, 6838, 3968}, '{-31917, 25976, -27740, -12591, -9068, 24437, 7152}}
    },
    '{
        '{'{19715, -8066, 22314, -23999, -10732, 804, 5444}, '{19408, -16272, 1967, -15734, 4333, -31384, 13278}, '{30555, -18901, -32705, 3999, -28780, 18886, 29961}, '{19900, 12891, -13713, 13731, 2387, -6324, -10990}, '{3441, -24758, 26850, -19231, 18347, -27005, -13428}, '{-25372, 3898, 20353, -18063, 23680, -11481, 29720}, '{-7494, -16092, -1693, 25413, 14470, 20483, -27422}},
        '{'{-9351, 4776, -1604, -19039, -8932, 23364, -28646}, '{-32032, -5896, 4461, -14413, -21303, -19019, 8389}, '{13217, 1671, 27261, 606, -14264, 12534, 23380}, '{25735, 18115, 26837, -16933, -24980, 19779, 6246}, '{-8364, -5817, -7597, 5343, -30464, -20859, 3419}, '{1131, -1122, -18487, -14381, 28167, 27797, 10213}, '{-8740, -19064, 18091, -22994, -24576, -25240, 691}},
        '{'{13862, 29785, -5046, -13837, -5406, -30085, -7849}, '{-17312, -25773, -3814, 23246, -26592, -5005, 6598}, '{-26783, 4524, 827, -22727, 23218, -22355, -2327}, '{-29564, 28089, -32675, 15707, -19055, 2467, 3778}, '{-32364, -27731, -6983, 13263, -32393, -16732, 20329}, '{-21826, -508, -15887, 24050, -9011, -23138, -2707}, '{-2217, 8930, -28253, 6729, -29478, 10167, 1562}}
    },
    '{
        '{'{30070, -3050, -7732, -1329, 32098, -4518, 19507}, '{-1050, 18222, -16688, 32317, 26044, 23343, 30714}, '{14440, -28032, -29302, -12341, 22413, 28999, -28066}, '{5638, 7853, 15605, -27234, 13839, 14505, 6310}, '{13621, -29781, -11694, -4729, -29476, 19265, 5801}, '{31554, 23666, -21668, 8526, -7451, -6949, -778}, '{-24476, 18847, -22307, 29874, 7676, -8018, -7587}},
        '{'{-24974, -12639, 4876, -12576, 9961, 9040, 25666}, '{-10808, -3085, -30595, -23414, -11664, -25894, -15205}, '{-7496, -9096, 28993, -13888, -30011, -20648, -8926}, '{-28721, -14333, 23228, 19694, -24923, 31915, 18131}, '{11096, 32326, -24940, -7290, 3868, -11661, 4998}, '{-27838, 16988, 24540, 3686, -7323, -12933, -12603}, '{-19347, 9545, -32668, 21174, -23731, -26731, 22011}},
        '{'{-7521, 20049, 19491, -7955, 15603, 14586, -1656}, '{23294, 9497, -16363, -9811, 17637, 6102, -7792}, '{-2919, 25582, -29577, 9893, 8063, 30081, 30085}, '{18118, 6540, -29350, -23990, -1029, 21430, 7246}, '{9022, 26184, -1849, 32557, -13179, 15919, 29371}, '{-11094, 20931, -26486, 21234, -31431, 3547, -19111}, '{-15997, -27523, -5426, -28846, -31547, 14010, -30844}}
    },
    '{
        '{'{23569, -23867, 8639, 16734, -23912, -12669, -3771}, '{-24152, 4260, 24122, 9393, -29257, -21864, -32095}, '{1938, 24417, 12750, -7439, -25465, 18357, -3349}, '{28718, 32240, -1036, 10879, -1119, 8529, 21661}, '{-4596, 28278, 10030, 27510, -3808, 7970, 16499}, '{-27049, -5508, -3687, -4946, -22030, 24427, -460}, '{24553, -19858, 5696, -29364, 28534, -21943, 4242}},
        '{'{19204, 18183, 2691, 9264, -5044, -26331, -20364}, '{9709, -22992, 6253, -22574, -22349, 10801, 11335}, '{16218, 11697, -12306, 5405, 20995, -24502, -428}, '{-9750, 11585, 6007, -29164, -29488, -27606, 5618}, '{16412, 1434, 2903, 3252, -26320, 14274, -6554}, '{-7415, -25342, -21132, 31596, -2327, 13145, 13692}, '{-7307, -32156, -28582, -7100, 25193, 9738, -12276}},
        '{'{22120, 10465, -5723, -12121, -23648, 25978, 11553}, '{-23654, -32669, 23769, -30414, 26968, 31954, 22292}, '{13022, 32412, -31160, 21778, -2663, -7272, -25049}, '{-21270, -18821, 16668, -2408, -20846, 32451, 14508}, '{16083, 26925, 11062, -16384, 26762, 21187, 30598}, '{5851, 14179, 10681, 28614, 19347, 25762, -30670}, '{14578, 4966, -30700, -25941, -19850, 26752, 5604}}
    },
    '{
        '{'{-9875, -20375, 7874, 24801, -8564, 1807, -13194}, '{-17887, -5993, 1932, 3973, -986, 28417, -32502}, '{11270, -131, -27386, 8806, -4186, 12619, 30066}, '{25941, -4738, -13966, -9550, -205, -4862, -25268}, '{4765, 22025, -23949, -7224, -28283, -9612, 24757}, '{2283, 20673, 32555, -1457, -21442, -5812, 14895}, '{-9652, -2411, 16504, -18670, 14681, -7667, 16606}},
        '{'{3676, 20716, -22423, -21291, 11782, 12900, -12752}, '{-6616, 9114, -25442, -25211, 14479, 13247, -21019}, '{11301, -453, -16783, -20385, 14688, 2544, 14544}, '{-26336, 62, -5750, 27020, -2467, -16576, -2659}, '{6490, -30745, -24426, 24979, -13947, 2852, -3501}, '{16511, 1508, 9989, -17060, 18892, 23706, 12017}, '{-7085, 12172, 2022, -7033, -13132, -32176, -9827}},
        '{'{-15360, -12585, -1329, 32586, 32508, 28291, 4669}, '{18755, -21360, -22672, 9673, 7764, 116, 25317}, '{7935, 824, 30014, 23480, -9680, -11119, 26485}, '{8121, 3593, 12780, 21694, -6065, 25318, 23758}, '{-7775, 26500, -5232, 2276, -30905, 23870, 16151}, '{32603, 26990, -24569, 6653, 8982, 1890, -5986}, '{26358, 1616, 25755, -16849, 20975, 626, -17909}}
    },
    '{
        '{'{22487, 22350, -20505, -7394, -30630, -1758, -5578}, '{-6319, -9565, 23623, 7021, 16187, -19856, 4517}, '{-3004, -24139, -5107, 22629, -3309, 32619, 11528}, '{-25760, -14639, -2875, -5764, -24476, -31359, 765}, '{-11107, -27771, -8240, 20710, 12792, -26712, -30058}, '{-13282, -18177, -9709, 9988, 21140, -25750, -13750}, '{123, 15811, -810, 6460, 27365, -2822, -14755}},
        '{'{-3415, -27096, 26812, -23343, -3405, 1320, 14395}, '{2538, -23074, 18973, 14561, 7774, 23790, 11941}, '{20862, 10456, -752, -25757, 23719, 7837, 25084}, '{-13247, -16617, 27848, 1408, 1111, 3877, -10897}, '{-5697, -5734, 21209, -19111, 15494, 14552, 17911}, '{27087, -7067, -15063, 26513, 32720, 3952, 3115}, '{-15250, 19909, 20854, -29805, -9489, 14102, 28013}},
        '{'{8075, 31243, -17503, -8313, -6025, -28390, -7632}, '{-21305, 12527, -13642, 21088, -28316, -6318, -26025}, '{9621, -27138, 18946, 11528, 23818, -5883, 3366}, '{-25690, -23964, -11839, 26229, 571, -12636, 17285}, '{18693, 6182, 11939, -10152, -16463, 5839, -684}, '{-9870, -23287, 12279, 7300, 31665, -13288, -22946}, '{19842, 24403, 20355, -12723, -31477, 24973, 2532}}
    },
    '{
        '{'{2129, -7014, -20538, 18095, -2462, 30229, -20588}, '{-26966, -24710, 18873, -15215, -3483, -12327, -4876}, '{6613, 16567, -16796, -4924, -28561, 21730, 19211}, '{12258, -26527, -14098, -1645, -16528, -11253, 7137}, '{13849, 5217, -27297, 18733, 19206, -17831, -20648}, '{-5651, -30170, 4147, 9232, 24471, 28378, 21251}, '{1882, 12718, -24966, 21917, -3326, -32123, 21881}},
        '{'{-28729, 23311, -9394, -23133, -10060, -10905, 16246}, '{-9977, 10931, -21146, -32007, -23629, -12387, 4791}, '{625, 8587, 27075, 5837, -20614, 3383, 32344}, '{-30213, -17156, 20984, -2236, 27765, -18061, -554}, '{-27463, -1699, 6758, -19573, 16078, -25006, 28633}, '{3308, -4093, 165, 1415, 18205, 9294, 28427}, '{-21559, 16907, -1264, -25540, 27259, 24679, 14015}},
        '{'{699, -10111, -18542, -20811, -19172, -15936, 29525}, '{-20776, -2487, 15240, -8238, -29301, -22052, -9867}, '{14259, 27473, -3657, -29681, -32637, 29802, 27096}, '{16597, 3356, -4294, -20779, -31154, 2927, -7359}, '{4940, -31477, -6887, -15001, 30475, 25434, -27923}, '{-10846, 30593, 19454, 17040, 11521, -22000, -30175}, '{19489, 23724, 1510, 9000, -5816, 26829, -31638}}
    },
    '{
        '{'{595, -27918, 17824, -11369, 16708, -27233, 8854}, '{-9152, 7909, 32031, 79, 24659, 23311, 11059}, '{32249, 11660, -5459, -27638, 22004, 9833, 9040}, '{-5050, 30741, 11998, -31037, 17744, -10944, 9345}, '{-6350, -17568, -16021, 29691, -28206, 18770, -23879}, '{-12906, 7951, -23665, 11804, -29369, -19173, -18216}, '{-28359, 19258, 10456, -2100, -14067, -26734, 16462}},
        '{'{-24626, 22292, -27065, -2377, -4820, -1813, -8971}, '{19547, -10196, -24817, 10237, -14761, -26677, 1613}, '{8702, -25187, -10657, -3986, -16686, 7812, -3556}, '{30401, -6095, -27727, -13993, 15929, 7888, -25559}, '{-23078, 18160, 9410, 7087, 18705, 31764, -1370}, '{-31424, 32390, -16148, -3434, 18511, 6218, -15198}, '{28328, 6822, 19446, -10603, -8414, 8565, 11424}},
        '{'{18858, -6785, 15660, -32157, 30505, -9479, 15207}, '{-28773, 14075, -30416, 21887, -14710, 13636, -23279}, '{-9469, 24165, 22110, 29143, -22243, -19866, 1659}, '{7326, -11061, -3646, 19933, -25284, -5497, 6835}, '{-26380, 10825, 11735, -18496, 30704, -3695, 13992}, '{-16141, 2581, -2466, 14234, 3215, 2800, 14097}, '{-9974, -14703, -18301, 19431, -439, -15587, -9021}}
    },
    '{
        '{'{27079, 4560, 2274, -20860, -7747, -2214, -7068}, '{14470, 28704, 11345, -14729, -30346, 18165, -26331}, '{14967, -15077, 29747, 13902, 16315, 5718, -31137}, '{-6136, -13000, -9443, -1380, 18399, 21922, -24390}, '{22399, -28802, -12335, -27172, 26735, -8560, -4152}, '{-10693, 12535, -31764, -11257, -5236, 13600, 20180}, '{-11541, 28747, -29475, -31704, -19456, 24788, 25709}},
        '{'{14940, -819, -19291, 31151, 29245, 4199, -2126}, '{25156, -24082, -25652, 16057, 9079, 12261, -28688}, '{-19324, -1431, 2596, 29008, -22062, 16549, -23842}, '{-16011, 26094, -8925, -10320, 13952, 22065, -13127}, '{20745, -10190, -5407, 9392, 24561, 29196, -4410}, '{15996, -13837, -18524, 13411, -3738, -11228, 23838}, '{22130, 23699, -4698, 29100, -16349, -11506, 22557}},
        '{'{16307, 16444, -19464, -25263, 23363, 26397, -20325}, '{15491, 17441, 32501, -11853, -28810, 1435, 3300}, '{-24520, -26347, -3417, -12566, 7498, -13795, -5903}, '{-5219, 957, 9786, -26856, -12174, 11536, -26176}, '{-12444, 30690, -17797, -6131, 769, 28411, -28414}, '{1858, 10387, -22028, -12550, -27188, -29026, 1575}, '{-555, 5709, 2993, 1306, 12659, 17548, -29455}}
    },
    '{
        '{'{17344, -22271, -12892, -16630, 20330, 22816, -23042}, '{-25316, 27322, 15042, 2780, 29761, 17613, 31059}, '{6703, -17839, -3676, -825, -6859, 9926, -11639}, '{19983, -9454, -31587, 29365, 3004, 12842, -30254}, '{23170, -21731, -18031, 18467, 31608, 3347, -12400}, '{-12777, -24948, 4451, -25747, 14008, 26306, -25836}, '{15491, -20399, -13396, -30682, 23594, -9270, -19931}},
        '{'{362, -28120, 18287, -20709, -18812, 1459, 27030}, '{10917, 6947, 542, 18183, -25640, 13912, -32529}, '{-18545, -5750, -25453, 2893, 6119, 22328, -26651}, '{16359, 10130, 7623, 16444, 24600, -20320, -29332}, '{-8921, -1164, 31848, 13694, 367, 4212, 26596}, '{-18454, 20496, -19532, -10022, -20504, 26832, 25390}, '{-25376, 2654, 18260, 20247, -12657, 20652, 14931}},
        '{'{-27529, -14793, -19102, -21093, -26323, 23522, -19119}, '{-28969, 32155, 28237, -32336, 26583, 11102, -10875}, '{-7815, 20711, -3359, 17265, -19486, 18204, -4876}, '{15425, -14268, -1323, -5688, -26884, -32398, 7073}, '{-19082, 7651, 26160, -11165, 8153, 13893, -18495}, '{18019, 26695, -5631, 16513, 4295, -20839, 9316}, '{-13747, 7788, 3250, -31333, -28576, 17963, -28909}}
    },
    '{
        '{'{-9886, -15059, -24476, -11952, 28784, 27882, 21369}, '{23467, 15811, 14856, 30931, 31662, -26048, -32396}, '{28564, -29600, -14878, -3221, -1659, -20139, -26344}, '{9218, -9731, 31741, 3527, 29804, 2251, 243}, '{-228, 16758, -19617, -28607, -30256, 22898, 28882}, '{11662, 15893, -2961, -10385, 6341, -23775, 15978}, '{-11134, 12827, 27368, -11913, 15507, -28785, 4935}},
        '{'{18412, 6941, 17827, -13599, -18128, -31823, -31920}, '{-3912, 16703, -25128, -6726, -19579, -2253, 21754}, '{21053, 19562, 27091, 23825, -30675, 5088, 9790}, '{19478, 29921, -8602, 28297, 31493, 17740, 30269}, '{-5974, -15625, -11888, 3387, 28945, 31940, 17724}, '{-26983, 5262, -31891, -24771, -3915, -32687, 28189}, '{2246, -20452, 16074, -379, 31204, -19996, 31060}},
        '{'{12215, -11790, -28494, -29098, -26443, -6390, -4565}, '{-21573, -6754, -26821, 9358, 26611, -19024, -11656}, '{30077, 1080, -11839, 1896, -121, 31685, 10383}, '{8823, 3049, -22220, 6432, 11351, 14286, -29790}, '{22045, -10189, 24025, 8629, -5372, -27456, 3963}, '{-14182, -6700, 2437, -1670, -25768, -30447, -22588}, '{-30408, -22368, -19215, -32431, -2488, 16457, -15644}}
    },
    '{
        '{'{-2657, 26974, -4791, 29036, 3248, -32029, -19040}, '{5390, -11715, -4777, 24992, 26936, -24164, -28501}, '{-19359, -16206, 27438, 26732, -10424, -13915, -5512}, '{10242, -23791, -12145, -15677, -23211, 22000, -3342}, '{-13219, -18587, 15480, -17770, -27438, -8697, 9015}, '{-22351, -11238, 29432, 25220, -17299, 24665, 29722}, '{-324, 10483, -12689, -10669, -17842, -28014, 11385}},
        '{'{19040, -22181, -5340, 32102, 32148, -6785, -27156}, '{24963, 18066, 8397, -6093, -3535, -481, -1567}, '{22162, 18700, -9617, 32731, 30951, -21662, -8377}, '{-4514, 6957, 3792, -22463, -14248, 14608, -26323}, '{22911, 6363, 165, -15950, 14744, 1968, 1228}, '{-23548, 21488, -11341, 1198, 31784, -4210, 11505}, '{-18038, -25189, 3406, -27802, 5517, 19972, -11562}},
        '{'{21775, 7197, -23602, -9046, 32409, -15157, 12767}, '{-8997, 18966, -25490, -3285, 1492, 3767, -17667}, '{17538, -8551, 26237, -1928, -14720, -12961, -32584}, '{7278, 11974, -27694, -1450, 10430, -257, 7726}, '{-19717, 5209, 19149, 18060, -26306, 16677, 20435}, '{14495, -27785, -24676, 26939, 30200, -3757, -4312}, '{9576, -2695, -8615, -20497, -28899, 31516, -7116}}
    },
    '{
        '{'{32042, -5494, 3796, -27375, 25216, 11943, 28710}, '{1506, -7999, -16848, -18218, -25555, 1146, 2737}, '{30230, -3865, -10754, -17060, -15039, -31403, 30530}, '{-18912, -13902, 25926, 27238, 23459, -6155, 25060}, '{-14185, -16397, -30598, 18514, 5222, -16295, 25326}, '{30799, -29583, -24421, 24405, 1537, 2313, -20365}, '{-30895, -20085, -11200, 2295, 5955, -12807, -835}},
        '{'{-8138, -15068, 31188, -4994, -24557, 1007, -12603}, '{4820, 23165, -16706, -828, 21673, 16592, -13680}, '{2233, -16763, -6048, 2326, -2941, -14968, 21310}, '{-6308, -31575, 10058, 24678, -22948, 15455, 18540}, '{-31861, 21410, 16475, 18225, 12871, 26023, 27494}, '{-17545, -966, 29701, 1097, 18264, 12428, 2792}, '{25825, 28475, -11570, 14317, 11791, -23548, 30614}},
        '{'{-31052, 14402, -12473, -25235, -5816, 3333, 25127}, '{-24241, 12111, -4311, 15321, 662, -17959, -23335}, '{-11373, 7998, -23779, 9993, 28043, -21635, -10141}, '{-486, -21657, -2817, 3794, -25016, -16129, 30337}, '{-8349, 6770, 6385, 32430, 9527, 26122, -16694}, '{5400, -1537, -10913, 29739, -3109, -31091, -11314}, '{20535, -26619, -7785, 22570, -27033, -17359, 17765}}
    }
};
