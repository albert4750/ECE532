localparam bit signed [0:46][15:0] Input1 = '{16'd28679, -16'd30103, -16'd13327, -16'd1911, 16'd6838, 16'd3968, -16'd31917, 16'd25976, -16'd27740, -16'd12591, -16'd9068, 16'd24437, 16'd7152, 16'd19715, -16'd8066, 16'd22314, -16'd23999, -16'd10732, 16'd804, 16'd5444, 16'd19408, -16'd16272, 16'd1967, -16'd15734, 16'd4333, -16'd31384, 16'd13278, 16'd30555, -16'd18901, -16'd32705, 16'd3999, -16'd28780, 16'd18886, 16'd29961, 16'd19900, 16'd12891, -16'd13713, 16'd13731, 16'd2387, -16'd6324, -16'd10990, 16'd3441, -16'd24758, 16'd26850, -16'd19231, 16'd18347, -16'd27005};
