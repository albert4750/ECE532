localparam bit signed [0:2][47:0] Bias3 = '{48'd5551, 48'd5363, 48'd5546};
