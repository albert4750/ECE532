logic signed [15:0] layer3_weight[3][12][3][3] = '{
    '{
        '{'{-25621, 26750, 4483}, '{28992, -475, 20983}, '{-14681, -11252, -21676}},
        '{'{3531, -18100, 5752}, '{-28302, -37, -11345}, '{4409, 18581, 28524}},
        '{'{524, 22511, 17041}, '{-9817, -24673, -22929}, '{-26979, 6583, 2497}},
        '{'{9509, -17920, -23785}, '{-27763, 136, -17964}, '{-18379, -30510, 31056}},
        '{'{12045, -18040, 11654}, '{-7781, -21339, 419}, '{-472, 28314, 6494}},
        '{'{-31796, -583, -14035}, '{-28848, -4806, 7319}, '{-13570, 23794, -32022}},
        '{'{-31800, 8183, -1034}, '{-13872, -4875, 11133}, '{-18926, -27702, -30833}},
        '{'{25062, -26755, -27816}, '{-2076, 22255, 19264}, '{-25213, 20442, 19348}},
        '{'{5103, 11439, 18878}, '{29025, 3096, 27346}, '{-2264, -18295, -19128}},
        '{'{27847, 32220, 6127}, '{16681, -2285, -9514}, '{9539, 30711, -26674}},
        '{'{11391, 28279, 8002}, '{-18729, -12053, -27624}, '{-12716, -10589, 30586}},
        '{'{19886, 4640, -19678}, '{22058, 860, 6181}, '{16612, -3246, -15305}}
    },
    '{
        '{'{-26774, -21981, -16409}, '{16739, 23617, 14685}, '{13972, -27419, 18787}},
        '{'{-19666, 7522, 91}, '{30782, 26686, -24079}, '{18683, -21938, 4970}},
        '{'{-18274, -17061, -20429}, '{-9724, 14020, 902}, '{16105, -215, 7427}},
        '{'{2727, -22036, 23652}, '{6555, 16013, 16684}, '{6400, -22710, -29987}},
        '{'{-31922, -31616, -13056}, '{-26528, 18292, -16629}, '{-10211, 23941, 18501}},
        '{'{-11591, -23266, -5358}, '{4714, -8176, -6281}, '{11601, 13515, -22519}},
        '{'{-14455, -9510, -7092}, '{26304, -27417, -6244}, '{-14602, 11085, 29527}},
        '{'{11194, 10873, 7600}, '{-4709, -22677, -3943}, '{-26668, -10129, -10676}},
        '{'{-14824, -12539, -19422}, '{-16308, 11451, -29141}, '{9167, -23749, 3349}},
        '{'{7652, -25103, 6654}, '{-26260, -14836, -21648}, '{31842, 25221, 16148}},
        '{'{-31108, -1377, 30562}, '{26903, -2541, -26027}, '{-29905, -30726, 20230}},
        '{'{68, -11063, 32280}, '{13231, -8288, 6090}, '{27354, -11813, 1296}}
    },
    '{
        '{'{-31006, -9066, -27523}, '{-15332, -20196, 2673}, '{24526, -25755, -21927}},
        '{'{-15227, 17986, -10845}, '{25291, 15283, 19021}, '{-10269, 27320, -8737}},
        '{'{21982, 23813, 26653}, '{22619, 30713, -16459}, '{29121, -2755, 20968}},
        '{'{19610, -25316, 999}, '{-13913, 15969, 105}, '{23215, -18323, -2144}},
        '{'{20857, -20220, 21942}, '{2432, -7925, 8371}, '{16995, -15420, -8422}},
        '{'{-497, -9743, -7460}, '{31594, 21392, 29556}, '{-7098, -5384, 26719}},
        '{'{17410, 12796, 32017}, '{-21262, 12097, 14496}, '{-30495, 9638, 2628}},
        '{'{-14498, -25340, -3077}, '{-14001, 21631, 20757}, '{-28807, 30067, 9318}},
        '{'{30474, -20208, -30718}, '{14126, 17085, 22702}, '{21614, -14048, 24807}},
        '{'{-18537, -28995, -7807}, '{-21212, 3929, 264}, '{22063, 27483, 17408}},
        '{'{-32605, 23578, -27458}, '{-26769, 2996, -16406}, '{9878, 23199, 3713}},
        '{'{-6307, 2307, -32509}, '{9570, -27532, 24740}, '{22954, -3730, 13332}}
    }
};
