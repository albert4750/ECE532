localparam bit signed [0:2][0:26][19:0] Input9 = '{
    '{20'd98, 20'd35, -20'd55, 20'd90, 20'd55, -20'd102, -20'd10, -20'd106, 20'd76, 20'd79, -20'd30, -20'd38, -20'd77, 20'd102, -20'd82, 20'd80, -20'd67, 20'd60, -20'd81, 20'd122, -20'd24, 20'd0, 20'd10, 20'd75, 20'd13, -20'd57, -20'd34},
    '{-20'd122, 20'd45, 20'd117, 20'd30, -20'd113, 20'd41, 20'd38, -20'd75, 20'd43, -20'd46, 20'd7, 20'd92, -20'd63, 20'd41, -20'd62, -20'd14, -20'd36, -20'd50, 20'd101, 20'd91, 20'd118, -20'd28, 20'd31, 20'd93, 20'd50, 20'd124, 20'd46},
    '{-20'd35, -20'd14, 20'd33, -20'd116, 20'd96, 20'd105, -20'd48, -20'd62, 20'd72, 20'd115, -20'd3, 20'd10, -20'd16, 20'd90, 20'd27, 20'd56, -20'd8, -20'd63, 20'd64, 20'd69, -20'd40, -20'd94, 20'd79, -20'd125, 20'd60, 20'd110, 20'd37}
};
