localparam bit signed [0:7][36:0] Bias2 = '{37'd91918, -37'd146106, 37'd8658, 37'd180660, -37'd102780, -37'd121131, -37'd160817, -37'd51809};
