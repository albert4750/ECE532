localparam bit signed [0:10][15:0] Output0 = '{16'd19185, -16'd24112, -16'd15503, -16'd6058, -16'd28847, 16'd21991, -16'd29028, -16'd8151, -16'd2454, 16'd5023, -16'd23576};
