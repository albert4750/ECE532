// constants
//
// Global constants.

`ifndef ECE532_CONSTANTS_SVH
`define ECE532_CONSTANTS_SVH

package constants;

    parameter int DSP_A_WIDTH = 25;
    parameter int DSP_B_WIDTH = 18;
    parameter int DSP_OUT_WIDTH = 48;

endpackage : constants

`endif  // ECE532_CONSTANTS_SVH
