localparam bit signed [0:2][47:0] Bias3 = '{48'd236097, 48'd2006738, 48'd368489};
