logic signed [15:0] layer2_weight[10][20][1][1] = '{
    '{
        '{'{-29293}},
        '{'{-26644}},
        '{'{19436}},
        '{'{14776}},
        '{'{3606}},
        '{'{16470}},
        '{'{-13844}},
        '{'{6373}},
        '{'{-9668}},
        '{'{23202}},
        '{'{-24003}},
        '{'{-7242}},
        '{'{1062}},
        '{'{-4395}},
        '{'{5084}},
        '{'{8880}},
        '{'{-28254}},
        '{'{-21571}},
        '{'{-22847}},
        '{'{-4938}}
    },
    '{
        '{'{27501}},
        '{'{-1810}},
        '{'{16529}},
        '{'{-26060}},
        '{'{10530}},
        '{'{12203}},
        '{'{8333}},
        '{'{-12271}},
        '{'{3871}},
        '{'{-14827}},
        '{'{-28446}},
        '{'{7789}},
        '{'{-4479}},
        '{'{-443}},
        '{'{-31825}},
        '{'{-17166}},
        '{'{-15194}},
        '{'{-4289}},
        '{'{1183}},
        '{'{-19620}}
    },
    '{
        '{'{-1946}},
        '{'{11002}},
        '{'{-3982}},
        '{'{-23312}},
        '{'{18244}},
        '{'{2469}},
        '{'{-16505}},
        '{'{-28093}},
        '{'{15414}},
        '{'{18453}},
        '{'{18581}},
        '{'{-21191}},
        '{'{13274}},
        '{'{-30398}},
        '{'{11996}},
        '{'{27439}},
        '{'{-7136}},
        '{'{4325}},
        '{'{26273}},
        '{'{25827}}
    },
    '{
        '{'{6074}},
        '{'{5024}},
        '{'{-22937}},
        '{'{29841}},
        '{'{-3191}},
        '{'{2659}},
        '{'{-2132}},
        '{'{6742}},
        '{'{6405}},
        '{'{-42}},
        '{'{20105}},
        '{'{-10122}},
        '{'{-28351}},
        '{'{-25923}},
        '{'{-28437}},
        '{'{4229}},
        '{'{-5910}},
        '{'{-28476}},
        '{'{10887}},
        '{'{-3146}}
    },
    '{
        '{'{19}},
        '{'{-22542}},
        '{'{11059}},
        '{'{2982}},
        '{'{-24587}},
        '{'{19191}},
        '{'{8845}},
        '{'{-8181}},
        '{'{-23721}},
        '{'{-27290}},
        '{'{-7626}},
        '{'{-17227}},
        '{'{-3509}},
        '{'{-30424}},
        '{'{30709}},
        '{'{29279}},
        '{'{-32253}},
        '{'{25079}},
        '{'{-8515}},
        '{'{17538}}
    },
    '{
        '{'{18375}},
        '{'{12546}},
        '{'{12569}},
        '{'{-12498}},
        '{'{-19067}},
        '{'{26640}},
        '{'{5234}},
        '{'{-3960}},
        '{'{17105}},
        '{'{-7048}},
        '{'{28018}},
        '{'{-12708}},
        '{'{-11698}},
        '{'{-12872}},
        '{'{-9722}},
        '{'{25165}},
        '{'{29240}},
        '{'{15324}},
        '{'{9987}},
        '{'{15852}}
    },
    '{
        '{'{-31429}},
        '{'{-4506}},
        '{'{18799}},
        '{'{-5116}},
        '{'{9216}},
        '{'{7883}},
        '{'{-15450}},
        '{'{19590}},
        '{'{18291}},
        '{'{-18796}},
        '{'{31224}},
        '{'{6854}},
        '{'{-112}},
        '{'{-27840}},
        '{'{16707}},
        '{'{27771}},
        '{'{19525}},
        '{'{8559}},
        '{'{-16323}},
        '{'{31015}}
    },
    '{
        '{'{-10949}},
        '{'{16592}},
        '{'{-24103}},
        '{'{25081}},
        '{'{-12322}},
        '{'{32027}},
        '{'{-9013}},
        '{'{23528}},
        '{'{-23616}},
        '{'{-11999}},
        '{'{1305}},
        '{'{4788}},
        '{'{16270}},
        '{'{-11600}},
        '{'{-22110}},
        '{'{22132}},
        '{'{5672}},
        '{'{-31822}},
        '{'{19134}},
        '{'{-910}}
    },
    '{
        '{'{-29397}},
        '{'{5751}},
        '{'{-2010}},
        '{'{10387}},
        '{'{7978}},
        '{'{23010}},
        '{'{-8474}},
        '{'{-11115}},
        '{'{24468}},
        '{'{-8870}},
        '{'{-11869}},
        '{'{8091}},
        '{'{-13693}},
        '{'{-13351}},
        '{'{-9348}},
        '{'{-3705}},
        '{'{-17148}},
        '{'{-15868}},
        '{'{30773}},
        '{'{-28279}}
    },
    '{
        '{'{-11324}},
        '{'{-9567}},
        '{'{2993}},
        '{'{11978}},
        '{'{-2153}},
        '{'{-17479}},
        '{'{31472}},
        '{'{-5152}},
        '{'{32589}},
        '{'{-21099}},
        '{'{-20388}},
        '{'{3095}},
        '{'{-3984}},
        '{'{-635}},
        '{'{-2115}},
        '{'{26626}},
        '{'{27904}},
        '{'{-14583}},
        '{'{5959}},
        '{'{8093}}
    }
};
