localparam bit signed [0:10][15:0] Output2 = '{16'd5038, -16'd16680, -16'd11195, -16'd14840, -16'd25603, 16'd14856, -16'd26667, -16'd2301, 16'd6584, -16'd11020, -16'd7843};
