localparam bit signed [0:63][47:0] Bias1 = '{-48'd73750, -48'd1936795, -48'd3083238, -48'd584210, -48'd4411302, -48'd2842454, 48'd4222716, -48'd1003057, -48'd1071679, 48'd2631557, 48'd500735, -48'd2115232, 48'd5195060, -48'd3913197, -48'd1499377, 48'd1346835, -48'd1638927, 48'd789306, 48'd2124514, -48'd4672087, 48'd7112176, -48'd1392247, -48'd3073184, -48'd2624254, -48'd3210454, 48'd2256575, 48'd4624432, -48'd5526184, -48'd3165883, 48'd1712140, -48'd2123610, -48'd4254706, -48'd936561, -48'd1972812, -48'd1560531, -48'd3015476, -48'd5603820, -48'd2893975, -48'd7507626, -48'd1109254, -48'd3747592, -48'd5791612, -48'd2463024, -48'd739067, -48'd1323010, 48'd4720413, -48'd33648, -48'd103537, -48'd1099709, -48'd1690, 48'd1693581, -48'd2174844, 48'd1329637, 48'd3866721, 48'd2587253, -48'd1474432, -48'd4136841, 48'd863252, -48'd10836764, 48'd2062876, -48'd3542350, -48'd4635987, -48'd844116, -48'd3990732};
