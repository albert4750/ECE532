logic signed [15:0] layer3_weight[3][10][5][5] = '{
    '{
        '{'{8341, -31280, 590, -14381, 24101}, '{20058, -23476, 13647, -19757, 3218}, '{19946, 30274, -3312, -21512, -16053}, '{-20509, 15881, 4473, 13641, -8418}, '{21526, -16790, 18708, 25193, 14803}},
        '{'{-19132, -21138, -27569, 21921, 27584}, '{-7313, 32655, 3405, -7287, -9167}, '{19178, 11402, 29041, 25191, -21982}, '{-18521, 14256, -15060, -8468, -7574}, '{22785, 10184, 21760, -6005, 2970}},
        '{'{-15906, -18581, -28758, -17645, -31915}, '{-8337, 26369, 9722, -23620, -7598}, '{3548, -25026, -20597, 23547, -9551}, '{7359, -3212, -15769, -8567, 25624}, '{22596, -13542, 20276, 3179, 27190}},
        '{'{-22059, -16690, -29539, -28799, 9422}, '{10496, 18959, -29279, -15712, -32003}, '{29427, -9499, -32571, -22626, 24054}, '{-5015, -19793, -6670, 7738, 32713}, '{-11915, -25721, 22526, 2974, 15701}},
        '{'{-7138, 22953, -9208, 30785, -12691}, '{19925, 27912, -21255, -3347, 21553}, '{4468, -1984, -30117, 14386, 19632}, '{-8743, 23197, 4679, 17946, 26079}, '{19854, -1159, 11027, 5246, -26488}},
        '{'{3111, -3171, -25321, -28851, -8152}, '{-21375, 857, 13784, 25374, 1449}, '{19280, 1404, 19262, 20299, -2201}, '{22343, 5734, 28117, -20520, 25893}, '{-17621, -26181, -20828, 8864, 23369}},
        '{'{17137, -7425, -10264, -29808, 28067}, '{-265, -20093, 5671, -15963, -10758}, '{23811, -21080, -17862, 19939, 32385}, '{-11773, -11765, 32131, 1134, 3582}, '{-1349, -2932, -18592, -6233, 6962}},
        '{'{-13568, -11722, -19402, 7791, 10071}, '{-7481, 1723, -12991, -15902, 14093}, '{-8264, -19426, -25259, -12719, 25239}, '{-29789, 9121, 25478, -22504, 21538}, '{31735, -18840, 12729, -32410, 4553}},
        '{'{-7528, 18141, 9733, 29936, 2992}, '{-29799, 5572, -10514, -26586, -1664}, '{32059, -30514, 19529, 14564, -4625}, '{6066, 16412, 17807, 29378, 3108}, '{-32121, 30673, -26977, -25429, 12329}},
        '{'{-2609, -29924, -20098, -24394, -6348}, '{-26506, 6826, 30456, 17823, -4010}, '{-1479, 23026, 11287, -19332, 4932}, '{-30144, 20369, -1850, -30652, -4917}, '{-10272, -11056, -4222, -4614, -1334}}
    },
    '{
        '{'{-29273, 25086, -25434, -10826, 7932}, '{1639, -27651, 9463, -12160, 31497}, '{-2485, -29268, -19404, 13521, -25244}, '{17769, 4783, -21819, 28137, 24112}, '{7590, -22492, -14972, -14597, -31759}},
        '{'{-18229, -25561, 4317, -11541, 28862}, '{-27987, 27083, -6358, 18592, -23679}, '{-27924, -15185, 3746, 27946, 21802}, '{29036, 7370, -24150, -28932, 14056}, '{28206, -23577, -8753, -17811, -12582}},
        '{'{18025, 1576, 10860, -3728, -18608}, '{-4693, 11100, 29120, -10689, 17452}, '{-13443, -1406, -20970, -8836, 6040}, '{-16468, -8365, -290, 6093, 21895}, '{11475, -1821, -20171, 501, -4802}},
        '{'{-2659, -7468, -29176, -19510, -15575}, '{-27742, 17582, 15293, 10955, -21251}, '{-7480, -18827, -31433, -16427, 18164}, '{6724, 303, 18951, 248, 28984}, '{-28587, -7082, -698, -32749, -4437}},
        '{'{13638, 30048, -29189, 20837, 17750}, '{18793, 7957, 26356, 23691, -2901}, '{-28605, 14048, 5021, -21611, -6959}, '{7493, -28945, -30245, -18175, -13663}, '{11688, -19093, -11161, -29959, 26283}},
        '{'{18483, 19429, 15710, 25042, -22090}, '{-6193, 28412, -28365, 18861, -23320}, '{-12963, 24708, 27320, -16976, -10376}, '{490, -1644, -31984, 1077, 2005}, '{17090, 21908, -4115, -23624, -11880}},
        '{'{7979, 32084, -7443, 14015, -7153}, '{-12959, -26344, 19800, -13976, 7771}, '{-8899, 29315, -22125, -7540, -28558}, '{-13012, 10058, 22921, 27327, 25564}, '{-11915, 16046, 9951, 32215, -16499}},
        '{'{-16827, -24915, 10216, 23687, 25897}, '{-7570, 400, -11086, -9433, -22493}, '{-30870, 14620, -6539, 9297, 10277}, '{-19967, 31185, 31006, 23586, 16244}, '{-19453, -16991, -30549, 27993, -14847}},
        '{'{-16030, -25160, 14129, -25497, -3288}, '{-5038, -7639, -24266, 23509, 18095}, '{-22948, -22657, -16447, -21719, 12070}, '{-10868, 18639, -27748, 13593, 6395}, '{-6926, 53, 24022, 24255, 7515}},
        '{'{9293, 1697, -5682, -22155, 9096}, '{-828, 18478, -29066, 4949, 16045}, '{7644, 30486, 16654, -22272, 20914}, '{-24091, -14154, 21682, 19337, -6367}, '{-21260, 9768, -23896, -25869, -6265}}
    },
    '{
        '{'{-31846, 3741, -6222, 12473, -6639}, '{638, -9974, 18731, -25666, 20705}, '{-63, 4838, 28541, -11501, -4899}, '{-11898, -25595, -13116, 17858, 32503}, '{-21080, 10728, 12240, -11449, -2136}},
        '{'{-21736, 17623, -10572, -29318, -9578}, '{-27095, -11514, 30840, 31950, -7629}, '{17063, -1025, 12824, 15391, 20116}, '{-16750, -3293, 15840, 23252, -27560}, '{23008, 5723, 16172, -8198, -31900}},
        '{'{-2606, -12138, 9698, -3169, -16718}, '{-8430, -5636, 3150, 3591, -32245}, '{-6465, 22218, 31673, -10950, 2598}, '{25769, -17450, -24640, -31710, 24785}, '{-3670, -8268, 11334, -21373, -1112}},
        '{'{-8325, 12379, 27596, -31065, -32555}, '{-11495, 32512, -20373, 12194, 1405}, '{31681, -26768, 2603, -30043, 12270}, '{-20373, 1497, 29655, -20694, -21005}, '{17092, -29004, -15929, -11171, 14337}},
        '{'{20503, -1833, -24232, 6489, -18107}, '{14230, 16369, -2992, -1697, 19696}, '{26304, -28174, 10179, 353, -4321}, '{-10810, 13364, 7744, 14088, -9448}, '{21574, -6837, 28612, 3902, 25845}},
        '{'{-31643, -20665, 26103, 17945, 27059}, '{-21718, -17787, 4005, 21380, 25340}, '{-26881, 11198, 10026, -1031, -29684}, '{-13552, -17223, -16827, -16371, -30965}, '{28630, -30358, -729, 5376, 16792}},
        '{'{-29840, -25957, 25463, -21858, 5336}, '{-9252, 9624, 5887, -21634, -19362}, '{2681, 14260, -24210, -25952, 24510}, '{24381, -2578, 17379, 11350, 15151}, '{4744, -16893, 8804, 23220, -26418}},
        '{'{-18628, -26908, -23749, 17873, -23621}, '{14291, -15016, -30632, 4195, 13554}, '{-20671, 24780, 22868, -17401, -31658}, '{-26836, 4856, 20687, 19488, 13345}, '{-29363, -6527, -4605, -24153, 8440}},
        '{'{17854, 8254, 20068, -25626, -5861}, '{21434, -27038, -31379, 20710, -12881}, '{-30823, 1360, 3312, 11378, -2561}, '{15561, 10905, 11712, 22287, 7669}, '{17488, -8470, -1539, 30308, 24583}},
        '{'{11671, -23311, -26328, -24026, 24429}, '{-13787, 9841, -6555, -6716, 11490}, '{20310, 4028, -29446, -21199, -3554}, '{3835, -2335, -2597, 19783, 16077}, '{26329, -31323, 18335, 21220, -6918}}
    }
};
