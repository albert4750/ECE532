localparam bit signed [0:7][36:0] Bias2 = '{37'd0, 37'd0, 37'd0, 37'd0, 37'd0, 37'd0, 37'd0, 37'd0};
