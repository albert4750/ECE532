localparam bit signed [0:146][7:0] Input2 = '{23, 125, 104, -76, -105, -6, -56, -87, 109, -68, -81, 15, -92, 65, -34, 101, -86, 126, -128, 83, 6, 93, -61, -97, -99, -112, 67, -102, 125, -122, 105, 101, -117, -47, -73, -3, -85, -61, -108, 91, 127, -9, 92, -114, -114, -48, 99, 63, -11, 102, -85, 27, -26, 87, 20, 123, -105, -94, -96, -63, -106, -107, 57, -60, -83, 104, 39, -104, -42, -111, 52, 90, 8, -123, 97, -42, 122, -46, -118, -66, -99, 11, 30, -57, -70, 94, -86, 85, -57, 25, 108, -74, -10, -45, -103, 45, -7, 106, 3, -12, 84, 113, -45, 121, -91, 33, 60, -20, 89, -121, 60, 37, -44, 122, -30, -112, 45, 104, 39, -95, -31, -63, 73, -41, -60, -104, -122, -31, -14, 127, -68, 88, -67, 116, 59, 119, -7, 74, -99, 111, 120, -100, 24, 3, 82, 21, -122};
