localparam bit signed [0:146][7:0] Input5 = '{-102, -111, 68, -85, 47, 94, -3, -36, 121, -56, 58, -101, -122, 7, 53, -9, 120, -102, -5, 75, -91, -35, 49, -108, 93, -9, 56, 61, 55, 92, 23, 57, 9, 0, -26, 19, 71, -78, -90, 67, 124, 30, -91, 56, -2, 105, 5, -69, 80, 90, 61, -97, 70, -39, 75, 17, -97, 31, -44, -38, -89, 117, 50, -54, -90, -60, -5, -89, -1, 79, -115, 35, 102, -5, 11, -25, -53, 112, -74, 36, -46, 75, 51, 34, 58, -48, -100, 9, -27, -120, 17, 112, 108, 92, 25, -34, -5, -27, 59, -5, 94, 121, -69, 58, -110, -116, 1, -101, -118, 67, 61, -112, -101, -4, -122, -128, -121, 25, -61, -69, 120, -12, 127, 36, 44, 85, -15, 118, 127, 72, -17, 38, 42, 97, 36, -60, -37, -115, 13, 41, -56, 6, -34, 12, -30, 3, 104};
