localparam bit signed [0:2][0:26][19:0] Input7 = '{
    '{-20'd99, 20'd33, -20'd13, -20'd75, -20'd9, 20'd51, -20'd42, 20'd118, -20'd121, -20'd23, 20'd113, 20'd9, 20'd54, 20'd0, -20'd45, -20'd8, 20'd36, 20'd81, 20'd20, -20'd11, 20'd112, -20'd125, -20'd2, -20'd86, -20'd63, -20'd108, -20'd92},
    '{-20'd60, 20'd80, -20'd16, 20'd47, 20'd10, 20'd109, -20'd24, 20'd94, -20'd37, -20'd85, -20'd65, 20'd31, 20'd20, 20'd70, -20'd119, 20'd60, -20'd37, -20'd17, 20'd35, -20'd45, -20'd52, -20'd110, -20'd15, -20'd54, 20'd98, 20'd97, 20'd43},
    '{20'd3, 20'd12, 20'd100, -20'd70, 20'd1, -20'd15, 20'd0, -20'd89, -20'd104, 20'd58, -20'd92, -20'd29, -20'd59, 20'd6, -20'd125, 20'd98, -20'd7, 20'd40, 20'd60, 20'd33, -20'd100, -20'd60, -20'd102, 20'd96, 20'd120, -20'd19, 20'd51}
};
