localparam bit signed [0:2][0:7][0:2][0:2][19:0] Weight3 = '{
    '{'{'{-20'd155543, 20'd224477, -20'd174986}, '{20'd28281, 20'd113122, 20'd0}, '{-20'd81307, 20'd51259, 20'd15908}}, '{'{-20'd21210, 20'd19443, -20'd76004}, '{-20'd91912, -20'd104285, 20'd10605}, '{20'd21210, 20'd31816, -20'd79539}}, '{'{-20'd17675, 20'd91912, 20'd68934}, '{20'd125495, 20'd54794, 20'd144938}, '{20'd106052, 20'd44188, 20'd42421}}, '{'{20'd125495, -20'd70701, -20'd90144}, '{-20'd144938, -20'd70701, -20'd26513}, '{-20'd40653, -20'd10605, -20'd45956}}, '{'{20'd97215, 20'd106052, 20'd21210}, '{20'd83074, 20'd1768, 20'd45956}, '{20'd61864, -20'd22978, -20'd30048}}, '{'{20'd47724, 20'd37118, -20'd37118}, '{-20'd21210, -20'd35351, 20'd35351}, '{-20'd49491, -20'd67166, 20'd30048}}, '{'{-20'd49491, -20'd60096, -20'd84842}, '{20'd14140, 20'd7070, -20'd44188}, '{20'd74237, 20'd81307, -20'd1768}}, '{'{-20'd37118, 20'd47724, 20'd84842}, '{20'd136100, 20'd53026, -20'd35351}, '{20'd7070, 20'd113122, -20'd1768}}},
    '{'{'{-20'd205474, 20'd207783, -20'd64644}, '{20'd293204, 20'd106200, 20'd2309}, '{-20'd161609, 20'd6926, -20'd85422}}, '{'{-20'd83113, -20'd87730, 20'd53100}, '{-20'd60026, -20'd62335, 20'd20778}, '{-20'd36939, 20'd27704, 20'd23087}}, '{'{-20'd46174, 20'd73878, -20'd25396}, '{-20'd64644, -20'd25396, 20'd18470}, '{20'd66952, 20'd106200, -20'd80804}}, '{'{20'd145448, 20'd50791, -20'd55409}, '{-20'd30013, -20'd32322, 20'd233178}, '{-20'd6926, -20'd66952, 20'd101583}}, '{'{20'd27704, -20'd2309, 20'd96965}, '{-20'd39248, -20'd30013, 20'd39248}, '{20'd73878, 20'd73878, -20'd6926}}, '{'{-20'd57717, 20'd110817, 20'd133904}, '{20'd55409, 20'd55409, 20'd53100}, '{-20'd62335, 20'd9235, 20'd217017}}, '{'{-20'd32322, -20'd80804, -20'd73878}, '{20'd41557, 20'd69261, 20'd76187}, '{20'd23087, -20'd13852, 20'd2309}}, '{'{-20'd13852, 20'd30013, 20'd133904}, '{20'd9235, -20'd39248, -20'd36939}, '{-20'd25396, 20'd87730, 20'd39248}}},
    '{'{'{-20'd125534, 20'd20542, -20'd141511}, '{-20'd269327, -20'd52496, -20'd100427}, '{-20'd223678, 20'd289869, -20'd205419}}, '{'{-20'd36519, -20'd20542, -20'd130099}, '{-20'd6847, -20'd102709, -20'd114121}, '{-20'd155205, -20'd9130, -20'd104992}}, '{'{20'd111839, 20'd18259, 20'd6847}, '{20'd114121, 20'd219113, 20'd102709}, '{-20'd11412, 20'd120969, -20'd9130}}, '{'{20'd15977, 20'd31954, 20'd15977}, '{20'd155205, 20'd66190, 20'd95862}, '{-20'd102709, 20'd13695, 20'd11412}}, '{'{-20'd43366, -20'd15977, 20'd11412}, '{20'd114121, 20'd95862, 20'd123251}, '{20'd127816, 20'd22824, 20'd45649}}, '{'{-20'd34236, -20'd70755, -20'd66190}, '{-20'd89015, -20'd98144, 20'd4565}, '{-20'd109557, 20'd29672, -20'd70755}}, '{'{-20'd2282, 20'd54778, -20'd79885}, '{-20'd38801, -20'd52496, -20'd38801}, '{20'd45649, -20'd2282, -20'd2282}}, '{'{20'd114121, 20'd15977, 20'd31954}, '{20'd38801, -20'd25107, 20'd100427}, '{-20'd27389, 20'd6847, 20'd98144}}}
};
