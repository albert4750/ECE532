localparam bit signed [0:46][15:0] Input0 = '{16'd9864, 16'd31757, 16'd18424, -16'd31865, -16'd2352, -16'd17416, 16'd31254, -16'd7688, -16'd8369, -16'd18471, -16'd26872, -16'd20765, -16'd24826, -16'd9007, 16'd9671, 16'd31188, 16'd5593, -16'd16446, -16'd2500, 16'd29072, 16'd19512, 16'd7026, 16'd3821, -16'd13673, -16'd24296, -16'd31740, 16'd2660, 16'd29676, -16'd30415, -16'd5801, -16'd10722, -16'd25034, -16'd8039, -16'd4332, -16'd8863, -16'd5787, -16'd21831, 16'd12695, -16'd613, -16'd31715, -16'd13407, -16'd10893, 16'd3893, -16'd30089, -16'd21581, -16'd27818, -16'd1546};
