localparam bit signed [0:146][7:0] Input7 = '{16, -33, -34, 126, 101, -90, 48, 60, -122, 112, 70, -9, -127, -17, 63, 65, -3, -107, -82, -128, 86, 36, 26, 20, -44, 103, -94, 113, -18, -67, 30, 27, 100, -55, -56, -76, -44, 23, -66, -80, 103, 59, -85, 42, 13, 120, -17, 121, -119, 27, -38, 101, -94, -58, 41, 109, -91, -122, -70, -43, -125, -53, 106, -117, 29, -50, 83, -102, -21, 127, -48, 35, -76, 17, -48, 10, 121, 60, 73, -29, 25, -1, 26, -77, -49, -101, 4, -26, 85, -25, 113, 53, -105, 108, 102, -21, -21, -106, -36, 110, -85, -122, 13, 77, 17, 40, -3, 94, 68, -110, 112, 2, -101, 8, 107, 79, -77, 87, 47, -65, 30, -115, -36, 46, 14, 114, 46, 45, -31, -124, -12, 10, -12, -65, -110, 100, 72, -9, -70, 73, 110, 13, -116, 29, -50, -24, -51};
