logic signed [7:0] output_weight[3][8][3][3] = '{
    '{
        '{'{-21, 16, 120}, '{126, 114, 37}, '{-114, 36, -14}},
        '{'{4, 114, -81}, '{0, -79, 37}, '{126, 75, -84}},
        '{'{-59, -24, 110}, '{-112, -112, -118}, '{-123, 23, 47}},
        '{'{-61, 38, 112}, '{-110, -34, 80}, '{-97, 42, -81}},
        '{'{-107, 97, -73}, '{-54, -20, -97}, '{-45, -62, 19}},
        '{'{31, -14, -109}, '{-89, 39, -67}, '{-31, 44, 116}},
        '{'{108, 54, 94}, '{-6, 103, 62}, '{76, 16, -48}},
        '{'{126, 6, 68}, '{-83, 84, 122}, '{30, -52, -5}}
    },
    '{
        '{'{53, 33, -38}, '{18, 6, -8}, '{2, 26, 110}},
        '{'{-103, -115, 63}, '{91, -66, -71}, '{-91, 45, 21}},
        '{'{-21, 120, -59}, '{121, -79, -103}, '{-116, -76, -58}},
        '{'{47, 125, -55}, '{10, -56, 90}, '{16, -33, -34}},
        '{'{126, 101, -90}, '{48, 60, -122}, '{112, 70, -9}},
        '{'{-127, -17, 63}, '{65, -3, -107}, '{-82, -128, 86}},
        '{'{36, 26, 20}, '{-44, 103, -94}, '{113, -18, -67}},
        '{'{30, 27, 100}, '{-55, -56, -76}, '{-44, 23, -66}}
    },
    '{
        '{'{-80, 103, 59}, '{-85, 42, 13}, '{120, -17, 121}},
        '{'{-119, 27, -38}, '{101, -94, -58}, '{41, 109, -91}},
        '{'{-122, -70, -43}, '{-125, -53, 106}, '{-117, 29, -50}},
        '{'{83, -102, -21}, '{127, -48, 35}, '{-76, 17, -48}},
        '{'{10, 121, 60}, '{73, -29, 25}, '{-1, 26, -77}},
        '{'{-49, -101, 4}, '{-26, 85, -25}, '{113, 53, -105}},
        '{'{108, 102, -21}, '{-21, -106, -36}, '{110, -85, -122}},
        '{'{13, 77, 17}, '{40, -3, 94}, '{68, -110, 112}}
    }
};
