localparam bit signed [0:31][47:0] Bias2 = '{48'd709, 48'd686, 48'd594, 48'd629, 48'd701, 48'd565, 48'd775, -48'd1045, 48'd763, 48'd753, 48'd803, 48'd904, 48'd882, 48'd782, 48'd850, 48'd541, 48'd450, 48'd562, -48'd468, 48'd717, 48'd905, 48'd702, 48'd270, 48'd611, 48'd675, 48'd843, 48'd971, 48'd384, 48'd587, 48'd556, 48'd601, 48'd899};
