localparam bit signed [0:7][33:0] Bias1 = '{34'd0, 34'd0, 34'd0, 34'd0, 34'd0, 34'd0, 34'd0, 34'd0};
