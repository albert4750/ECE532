localparam bit signed [0:7][47:0] Bias1 = '{-48'd248782, 48'd13796, 48'd12289, -48'd203021, -48'd448166, 48'd303605, 48'd8747, 48'd179097};
