localparam bit signed [0:46][15:0] Input5 = '{16'd13621, -16'd29781, -16'd11694, -16'd4729, -16'd29476, 16'd19265, 16'd5801, 16'd31554, 16'd23666, -16'd21668, 16'd8526, -16'd7451, -16'd6949, -16'd778, -16'd24476, 16'd18847, -16'd22307, 16'd29874, 16'd7676, -16'd8018, -16'd7587, -16'd24974, -16'd12639, 16'd4876, -16'd12576, 16'd9961, 16'd9040, 16'd25666, -16'd10808, -16'd3085, -16'd30595, -16'd23414, -16'd11664, -16'd25894, -16'd15205, -16'd7496, -16'd9096, 16'd28993, -16'd13888, -16'd30011, -16'd20648, -16'd8926, -16'd28721, -16'd14333, 16'd23228, 16'd19694, -16'd24923};
