localparam bit signed [0:46][15:0] Input7 = '{-16'd23990, -16'd1029, 16'd21430, 16'd7246, 16'd9022, 16'd26184, -16'd1849, 16'd32557, -16'd13179, 16'd15919, 16'd29371, -16'd11094, 16'd20931, -16'd26486, 16'd21234, -16'd31431, 16'd3547, -16'd19111, -16'd15997, -16'd27523, -16'd5426, -16'd28846, -16'd31547, 16'd14010, -16'd30844, 16'd23569, -16'd23867, 16'd8639, 16'd16734, -16'd23912, -16'd12669, -16'd3771, -16'd24152, 16'd4260, 16'd24122, 16'd9393, -16'd29257, -16'd21864, -16'd32095, 16'd1938, 16'd24417, 16'd12750, -16'd7439, -16'd25465, 16'd18357, -16'd3349, 16'd28718};
