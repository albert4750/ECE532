localparam bit signed [0:31][0:63][0:0][0:0][24:0] Weight2 = '{
    '{'{'{25'd2915205}}, '{'{-25'd1340994}}, '{'{-25'd116608}}, '{'{25'd174912}}, '{'{-25'd1107778}}, '{'{-25'd874562}}, '{'{25'd58304}}, '{'{-25'd1166082}}, '{'{25'd1924035}}, '{'{25'd2390468}}, '{'{25'd408129}}, '{'{-25'd4022983}}, '{'{-25'd2215556}}, '{'{-25'd1574211}}, '{'{-25'd1457603}}, '{'{25'd3381638}}, '{'{25'd932866}}, '{'{25'd1749123}}, '{'{25'd1107778}}, '{'{25'd2332164}}, '{'{-25'd1224386}}, '{'{-25'd1340994}}, '{'{-25'd1749123}}, '{'{25'd3556550}}, '{'{25'd1690819}}, '{'{-25'd1574211}}, '{'{25'd524737}}, '{'{25'd1340994}}, '{'{25'd116608}}, '{'{25'd757953}}, '{'{-25'd58304}}, '{'{25'd641345}}, '{'{25'd1515907}}, '{'{25'd1515907}}, '{'{25'd4081287}}, '{'{25'd1457603}}, '{'{-25'd2273860}}, '{'{-25'd1457603}}, '{'{25'd3265030}}, '{'{-25'd1340994}}, '{'{25'd4022983}}, '{'{25'd2973509}}, '{'{25'd1049474}}, '{'{-25'd1399298}}, '{'{25'd1282690}}, '{'{25'd1340994}}, '{'{25'd0}}, '{'{25'd1457603}}, '{'{-25'd408129}}, '{'{25'd1166082}}, '{'{-25'd349825}}, '{'{-25'd1982339}}, '{'{-25'd1340994}}, '{'{-25'd2040644}}, '{'{25'd3265030}}, '{'{25'd1107778}}, '{'{25'd58304}}, '{'{25'd1690819}}, '{'{-25'd1807427}}, '{'{25'd7404621}}, '{'{25'd1574211}}, '{'{-25'd3906375}}, '{'{-25'd6471755}}, '{'{25'd1924035}}},
    '{'{'{-25'd1824725}}, '{'{25'd1190038}}, '{'{-25'd793359}}, '{'{25'd714023}}, '{'{25'd1428046}}, '{'{-25'd1031366}}, '{'{25'd1745389}}, '{'{25'd1666053}}, '{'{25'd714023}}, '{'{25'd1586718}}, '{'{-25'd1269374}}, '{'{-25'd158672}}, '{'{25'd2618084}}, '{'{25'd1031366}}, '{'{-25'd2300740}}, '{'{25'd1666053}}, '{'{-25'd238008}}, '{'{25'd555351}}, '{'{25'd1110702}}, '{'{25'd317344}}, '{'{-25'd1269374}}, '{'{25'd5156832}}, '{'{-25'd872695}}, '{'{-25'd3173435}}, '{'{-25'd158672}}, '{'{-25'd555351}}, '{'{-25'd158672}}, '{'{-25'd158672}}, '{'{-25'd793359}}, '{'{-25'd2142069}}, '{'{-25'd476015}}, '{'{25'd1190038}}, '{'{25'd1269374}}, '{'{25'd158672}}, '{'{-25'd872695}}, '{'{-25'd1031366}}, '{'{-25'd952031}}, '{'{25'd396679}}, '{'{25'd1190038}}, '{'{-25'd952031}}, '{'{25'd0}}, '{'{25'd5474175}}, '{'{-25'd1586718}}, '{'{-25'd634687}}, '{'{25'd1904061}}, '{'{-25'd317344}}, '{'{-25'd2062733}}, '{'{-25'd1904061}}, '{'{25'd7774916}}, '{'{25'd2062733}}, '{'{-25'd872695}}, '{'{-25'd872695}}, '{'{-25'd2062733}}, '{'{25'd1190038}}, '{'{25'd10075656}}, '{'{-25'd714023}}, '{'{25'd1983397}}, '{'{25'd1507382}}, '{'{25'd2221405}}, '{'{-25'd1586718}}, '{'{-25'd1824725}}, '{'{25'd2618084}}, '{'{-25'd2142069}}, '{'{-25'd1031366}}},
    '{'{'{-25'd1044216}}, '{'{25'd1193390}}, '{'{25'd497246}}, '{'{25'd895042}}, '{'{25'd1740360}}, '{'{-25'd447521}}, '{'{25'd298347}}, '{'{25'd1193390}}, '{'{25'd2237606}}, '{'{-25'd2187881}}, '{'{25'd2734851}}, '{'{25'd944767}}, '{'{-25'd1640911}}, '{'{-25'd1790085}}, '{'{-25'd1790085}}, '{'{25'd2983474}}, '{'{25'd1889534}}, '{'{25'd298347}}, '{'{-25'd1143665}}, '{'{-25'd1243114}}, '{'{25'd646419}}, '{'{-25'd3132648}}, '{'{25'd2486229}}, '{'{25'd1093941}}, '{'{25'd149174}}, '{'{25'd1839809}}, '{'{25'd1988983}}, '{'{25'd3132648}}, '{'{25'd4624385}}, '{'{-25'd397797}}, '{'{25'd745869}}, '{'{-25'd1640911}}, '{'{-25'd198898}}, '{'{25'd1093941}}, '{'{25'd1342563}}, '{'{-25'd2237606}}, '{'{-25'd99449}}, '{'{-25'd497246}}, '{'{25'd596695}}, '{'{25'd1939258}}, '{'{25'd795593}}, '{'{25'd497246}}, '{'{25'd1243114}}, '{'{25'd1342563}}, '{'{-25'd1889534}}, '{'{25'd1342563}}, '{'{25'd1193390}}, '{'{-25'd1889534}}, '{'{-25'd2585678}}, '{'{-25'd248623}}, '{'{25'd1939258}}, '{'{25'd1243114}}, '{'{25'd1740360}}, '{'{-25'd696144}}, '{'{-25'd2038707}}, '{'{25'd1292839}}, '{'{-25'd2237606}}, '{'{25'd845318}}, '{'{25'd149174}}, '{'{25'd6315020}}, '{'{25'd99449}}, '{'{-25'd1988983}}, '{'{25'd1193390}}, '{'{-25'd2436504}}},
    '{'{'{25'd1963166}}, '{'{-25'd1243339}}, '{'{25'd2028605}}, '{'{25'd1308777}}, '{'{25'd1701411}}, '{'{25'd654389}}, '{'{25'd2682994}}, '{'{-25'd1505094}}, '{'{-25'd392633}}, '{'{25'd2094044}}, '{'{25'd1766849}}, '{'{-25'd458072}}, '{'{-25'd2224922}}, '{'{25'd1832288}}, '{'{-25'd1701411}}, '{'{25'd392633}}, '{'{-25'd196317}}, '{'{25'd1243339}}, '{'{-25'd3075627}}, '{'{25'd1897727}}, '{'{25'd130878}}, '{'{-25'd1505094}}, '{'{25'd392633}}, '{'{25'd916144}}, '{'{25'd2094044}}, '{'{-25'd719828}}, '{'{-25'd850705}}, '{'{-25'd1308777}}, '{'{-25'd4384404}}, '{'{-25'd719828}}, '{'{25'd785266}}, '{'{25'd65439}}, '{'{25'd1374216}}, '{'{25'd1505094}}, '{'{-25'd2028605}}, '{'{25'd1047022}}, '{'{-25'd1308777}}, '{'{25'd1635972}}, '{'{-25'd261755}}, '{'{25'd1112461}}, '{'{25'd2028605}}, '{'{-25'd2486677}}, '{'{-25'd327194}}, '{'{25'd65439}}, '{'{25'd458072}}, '{'{-25'd196317}}, '{'{25'd1374216}}, '{'{25'd130878}}, '{'{-25'd130878}}, '{'{25'd785266}}, '{'{25'd2486677}}, '{'{25'd261755}}, '{'{25'd2355799}}, '{'{25'd1308777}}, '{'{-25'd1243339}}, '{'{25'd2224922}}, '{'{-25'd588950}}, '{'{-25'd130878}}, '{'{-25'd1701411}}, '{'{-25'd8376175}}, '{'{25'd65439}}, '{'{-25'd2748433}}, '{'{-25'd1047022}}, '{'{25'd196317}}},
    '{'{'{-25'd668538}}, '{'{25'd1568492}}, '{'{25'd719964}}, '{'{-25'd1671344}}, '{'{25'd745676}}, '{'{-25'd257130}}, '{'{25'd874241}}, '{'{25'd437121}}, '{'{25'd1568492}}, '{'{-25'd179991}}, '{'{-25'd1105658}}, '{'{-25'd771389}}, '{'{-25'd2905567}}, '{'{25'd1439927}}, '{'{-25'd1902761}}, '{'{-25'd334269}}, '{'{-25'd1234223}}, '{'{-25'd2057039}}, '{'{-25'd77139}}, '{'{-25'd642825}}, '{'{25'd128565}}, '{'{25'd771389}}, '{'{25'd2211316}}, '{'{-25'd1619918}}, '{'{25'd1645631}}, '{'{25'd1774196}}, '{'{25'd745676}}, '{'{25'd0}}, '{'{-25'd617112}}, '{'{-25'd694251}}, '{'{-25'd899954}}, '{'{25'd1157084}}, '{'{-25'd1722770}}, '{'{25'd2314168}}, '{'{-25'd1388501}}, '{'{25'd1851335}}, '{'{-25'd1774196}}, '{'{25'd437121}}, '{'{-25'd1465640}}, '{'{25'd1388501}}, '{'{-25'd1697057}}, '{'{25'd1851335}}, '{'{-25'd2005613}}, '{'{25'd1105658}}, '{'{25'd1825622}}, '{'{-25'd797102}}, '{'{-25'd231417}}, '{'{-25'd2005613}}, '{'{25'd282843}}, '{'{25'd2108465}}, '{'{-25'd1619918}}, '{'{25'd1568492}}, '{'{25'd1568492}}, '{'{-25'd2854141}}, '{'{25'd1337075}}, '{'{25'd2262742}}, '{'{25'd308556}}, '{'{25'd2185603}}, '{'{25'd2237029}}, '{'{-25'd2956993}}, '{'{-25'd2725576}}, '{'{25'd257130}}, '{'{-25'd3265549}}, '{'{25'd565686}}},
    '{'{'{25'd1566521}}, '{'{-25'd734307}}, '{'{25'd3035134}}, '{'{-25'd2153966}}, '{'{-25'd1566521}}, '{'{25'd538492}}, '{'{-25'd636399}}, '{'{-25'd244769}}, '{'{25'd1615475}}, '{'{-25'd1713382}}, '{'{25'd1468613}}, '{'{25'd391630}}, '{'{-25'd538492}}, '{'{-25'd1419660}}, '{'{-25'd391630}}, '{'{-25'd2007105}}, '{'{25'd3084088}}, '{'{25'd342676}}, '{'{-25'd1419660}}, '{'{25'd489538}}, '{'{25'd342676}}, '{'{-25'd489538}}, '{'{-25'd979076}}, '{'{25'd6217130}}, '{'{25'd1517567}}, '{'{25'd1615475}}, '{'{25'd2056059}}, '{'{25'd3475718}}, '{'{25'd2692458}}, '{'{25'd587445}}, '{'{25'd1272798}}, '{'{25'd538492}}, '{'{25'd1174891}}, '{'{25'd342676}}, '{'{25'd1125937}}, '{'{-25'd1664428}}, '{'{-25'd1713382}}, '{'{25'd97908}}, '{'{-25'd1517567}}, '{'{25'd1615475}}, '{'{25'd1762336}}, '{'{25'd0}}, '{'{-25'd1664428}}, '{'{25'd146861}}, '{'{-25'd1076983}}, '{'{-25'd1958151}}, '{'{-25'd2398735}}, '{'{25'd3035134}}, '{'{-25'd1468613}}, '{'{-25'd391630}}, '{'{-25'd734307}}, '{'{25'd1566521}}, '{'{-25'd2007105}}, '{'{25'd2056059}}, '{'{25'd2202920}}, '{'{25'd48954}}, '{'{-25'd734307}}, '{'{-25'd1762336}}, '{'{-25'd342676}}, '{'{25'd4601655}}, '{'{25'd1909197}}, '{'{25'd244769}}, '{'{-25'd1125937}}, '{'{25'd2056059}}},
    '{'{'{-25'd525240}}, '{'{-25'd678434}}, '{'{25'd2166613}}, '{'{-25'd2735623}}, '{'{25'd459585}}, '{'{25'd2079073}}, '{'{-25'd525240}}, '{'{25'd1488179}}, '{'{-25'd1313099}}, '{'{-25'd2013418}}, '{'{-25'd2144728}}, '{'{-25'd1728913}}, '{'{-25'd2188498}}, '{'{25'd2451118}}, '{'{25'd43770}}, '{'{-25'd2626198}}, '{'{-25'd1597604}}, '{'{-25'd2210383}}, '{'{25'd569009}}, '{'{-25'd459585}}, '{'{25'd1597604}}, '{'{-25'd1072364}}, '{'{25'd196965}}, '{'{25'd1991533}}, '{'{-25'd153195}}, '{'{25'd1334984}}, '{'{-25'd2035303}}, '{'{-25'd1663259}}, '{'{25'd1203674}}, '{'{25'd787859}}, '{'{25'd1772683}}, '{'{25'd2035303}}, '{'{25'd1947763}}, '{'{25'd2013418}}, '{'{-25'd1116134}}, '{'{25'd2516773}}, '{'{-25'd65655}}, '{'{25'd2144728}}, '{'{-25'd1597604}}, '{'{25'd590894}}, '{'{25'd656549}}, '{'{-25'd612779}}, '{'{-25'd612779}}, '{'{-25'd2210383}}, '{'{25'd1882108}}, '{'{-25'd1181789}}, '{'{25'd2363578}}, '{'{25'd962939}}, '{'{25'd1159904}}, '{'{25'd1903993}}, '{'{25'd306390}}, '{'{-25'd984824}}, '{'{-25'd1947763}}, '{'{-25'd393930}}, '{'{-25'd2779393}}, '{'{25'd787859}}, '{'{25'd1072364}}, '{'{25'd393930}}, '{'{-25'd2079073}}, '{'{25'd1991533}}, '{'{25'd1072364}}, '{'{-25'd1488179}}, '{'{25'd1006709}}, '{'{25'd2166613}}},
    '{'{'{25'd350275}}, '{'{-25'd437844}}, '{'{25'd3721674}}, '{'{25'd1182179}}, '{'{-25'd1182179}}, '{'{-25'd1751376}}, '{'{25'd1576238}}, '{'{25'd481628}}, '{'{-25'd2320573}}, '{'{-25'd2233004}}, '{'{25'd2014082}}, '{'{25'd1488670}}, '{'{25'd218922}}, '{'{25'd744335}}, '{'{-25'd2364358}}, '{'{-25'd1357316}}, '{'{25'd525413}}, '{'{25'd2145436}}, '{'{25'd1313532}}, '{'{25'd262706}}, '{'{-25'd2320573}}, '{'{-25'd3196261}}, '{'{-25'd2583280}}, '{'{25'd2627064}}, '{'{25'd1751376}}, '{'{25'd306491}}, '{'{-25'd175138}}, '{'{25'd5560619}}, '{'{25'd2845986}}, '{'{25'd1926514}}, '{'{-25'd1707592}}, '{'{25'd306491}}, '{'{25'd2933555}}, '{'{-25'd1401101}}, '{'{-25'd3984380}}, '{'{-25'd1663807}}, '{'{-25'd1444885}}, '{'{-25'd1313532}}, '{'{25'd525413}}, '{'{25'd1225963}}, '{'{-25'd1313532}}, '{'{-25'd131353}}, '{'{25'd1138394}}, '{'{25'd2233004}}, '{'{25'd2233004}}, '{'{25'd656766}}, '{'{-25'd2627064}}, '{'{25'd5035206}}, '{'{-25'd1926514}}, '{'{25'd1313532}}, '{'{25'd1970298}}, '{'{-25'd2145436}}, '{'{25'd481628}}, '{'{25'd1094610}}, '{'{-25'd481628}}, '{'{-25'd394060}}, '{'{25'd919472}}, '{'{-25'd1620023}}, '{'{-25'd2320573}}, '{'{25'd5516834}}, '{'{25'd3240046}}, '{'{-25'd1970298}}, '{'{-25'd1357316}}, '{'{25'd1926514}}},
    '{'{'{25'd1611340}}, '{'{25'd867645}}, '{'{25'd3346630}}, '{'{-25'd1673315}}, '{'{25'd1735290}}, '{'{-25'd1983188}}, '{'{-25'd2107137}}, '{'{-25'd2355036}}, '{'{25'd805670}}, '{'{-25'd185924}}, '{'{25'd557772}}, '{'{25'd991594}}, '{'{-25'd2726884}}, '{'{-25'd929619}}, '{'{25'd1177518}}, '{'{25'd1611340}}, '{'{25'd1363442}}, '{'{25'd247899}}, '{'{-25'd5019945}}, '{'{-25'd1735290}}, '{'{25'd495797}}, '{'{-25'd1301467}}, '{'{25'd1859239}}, '{'{25'd1611340}}, '{'{-25'd61975}}, '{'{25'd929619}}, '{'{25'd2107137}}, '{'{-25'd2726884}}, '{'{25'd2850833}}, '{'{-25'd1673315}}, '{'{25'd2045163}}, '{'{-25'd495797}}, '{'{25'd1673315}}, '{'{25'd743696}}, '{'{-25'd185924}}, '{'{-25'd247899}}, '{'{25'd123949}}, '{'{25'd2169112}}, '{'{-25'd1363442}}, '{'{-25'd2293061}}, '{'{25'd1487391}}, '{'{25'd3904402}}, '{'{25'd2478985}}, '{'{-25'd61975}}, '{'{-25'd2169112}}, '{'{25'd0}}, '{'{25'd805670}}, '{'{-25'd2355036}}, '{'{-25'd1425416}}, '{'{-25'd309873}}, '{'{25'd1611340}}, '{'{-25'd247899}}, '{'{-25'd743696}}, '{'{25'd2355036}}, '{'{25'd7870778}}, '{'{-25'd929619}}, '{'{-25'd681721}}, '{'{-25'd2355036}}, '{'{25'd743696}}, '{'{25'd6259437}}, '{'{25'd247899}}, '{'{25'd2045163}}, '{'{25'd991594}}, '{'{-25'd1487391}}},
    '{'{'{-25'd1079215}}, '{'{-25'd503634}}, '{'{-25'd503634}}, '{'{-25'd359738}}, '{'{-25'd791425}}, '{'{-25'd2014536}}, '{'{25'd719477}}, '{'{-25'd2014536}}, '{'{-25'd2374274}}, '{'{25'd791425}}, '{'{-25'd863372}}, '{'{-25'd2446222}}, '{'{25'd8130090}}, '{'{25'd71948}}, '{'{-25'd1726745}}, '{'{25'd2302326}}, '{'{25'd2158431}}, '{'{25'd1510902}}, '{'{25'd4964391}}, '{'{-25'd719477}}, '{'{25'd2014536}}, '{'{25'd7698404}}, '{'{-25'd791425}}, '{'{-25'd3741280}}, '{'{-25'd647529}}, '{'{-25'd71948}}, '{'{25'd2230379}}, '{'{-25'd791425}}, '{'{25'd1798692}}, '{'{25'd2302326}}, '{'{-25'd2662065}}, '{'{25'd4316862}}, '{'{-25'd503634}}, '{'{25'd1438954}}, '{'{25'd5539973}}, '{'{-25'd2446222}}, '{'{25'd9137358}}, '{'{25'd2374274}}, '{'{-25'd71948}}, '{'{-25'd1942588}}, '{'{-25'd647529}}, '{'{25'd0}}, '{'{-25'd215843}}, '{'{25'd1007268}}, '{'{25'd71948}}, '{'{25'd4101019}}, '{'{-25'd1798692}}, '{'{-25'd1510902}}, '{'{25'd3813228}}, '{'{25'd1798692}}, '{'{25'd0}}, '{'{-25'd1582849}}, '{'{25'd791425}}, '{'{25'd1223111}}, '{'{25'd5324130}}, '{'{25'd935320}}, '{'{25'd863372}}, '{'{-25'd1079215}}, '{'{25'd791425}}, '{'{25'd935320}}, '{'{-25'd1367006}}, '{'{25'd1870640}}, '{'{25'd71948}}, '{'{25'd0}}},
    '{'{'{25'd1899682}}, '{'{-25'd523101}}, '{'{-25'd330379}}, '{'{25'd27532}}, '{'{-25'd688291}}, '{'{25'd1293986}}, '{'{25'd3496516}}, '{'{-25'd963607}}, '{'{25'd2119935}}, '{'{-25'd1046202}}, '{'{25'd495569}}, '{'{25'd2367720}}, '{'{25'd825949}}, '{'{25'd825949}}, '{'{25'd1321518}}, '{'{25'd3083542}}, '{'{25'd1459176}}, '{'{25'd495569}}, '{'{25'd1018670}}, '{'{25'd1376581}}, '{'{-25'd1046202}}, '{'{-25'd2587973}}, '{'{-25'd1404113}}, '{'{25'd468038}}, '{'{25'd1431644}}, '{'{-25'd2532909}}, '{'{25'd2147467}}, '{'{-25'd3468984}}, '{'{-25'd715822}}, '{'{25'd1486708}}, '{'{-25'd1349050}}, '{'{25'd468038}}, '{'{25'd881012}}, '{'{25'd82595}}, '{'{25'd1459176}}, '{'{-25'd1404113}}, '{'{-25'd1899682}}, '{'{-25'd578164}}, '{'{25'd2477846}}, '{'{-25'd1376581}}, '{'{-25'd1183860}}, '{'{25'd1734492}}, '{'{25'd2257593}}, '{'{25'd1183860}}, '{'{25'd1651897}}, '{'{-25'd1404113}}, '{'{25'd55063}}, '{'{25'd330379}}, '{'{-25'd165190}}, '{'{-25'd1817087}}, '{'{25'd110126}}, '{'{-25'd137658}}, '{'{25'd908544}}, '{'{-25'd220253}}, '{'{25'd715822}}, '{'{-25'd2395251}}, '{'{-25'd1624366}}, '{'{25'd1349050}}, '{'{25'd1844619}}, '{'{-25'd1899682}}, '{'{-25'd2505378}}, '{'{25'd220253}}, '{'{-25'd2367720}}, '{'{25'd1872150}}},
    '{'{'{25'd1512657}}, '{'{25'd126055}}, '{'{25'd2479077}}, '{'{-25'd1554675}}, '{'{-25'd336146}}, '{'{25'd840365}}, '{'{-25'd1176511}}, '{'{-25'd210091}}, '{'{-25'd1932840}}, '{'{25'd840365}}, '{'{-25'd210091}}, '{'{-25'd630274}}, '{'{25'd1134493}}, '{'{25'd2184949}}, '{'{25'd1302566}}, '{'{25'd2437059}}, '{'{-25'd2268986}}, '{'{25'd2100913}}, '{'{25'd1344584}}, '{'{25'd1386602}}, '{'{25'd378164}}, '{'{-25'd1134493}}, '{'{-25'd840365}}, '{'{-25'd1176511}}, '{'{25'd1344584}}, '{'{-25'd168073}}, '{'{25'd2142931}}, '{'{-25'd882383}}, '{'{25'd2479077}}, '{'{25'd42018}}, '{'{25'd672292}}, '{'{-25'd882383}}, '{'{-25'd840365}}, '{'{-25'd1218529}}, '{'{25'd1386602}}, '{'{25'd2268986}}, '{'{25'd1638712}}, '{'{25'd1134493}}, '{'{-25'd546237}}, '{'{-25'd336146}}, '{'{-25'd1260548}}, '{'{-25'd1638712}}, '{'{-25'd924402}}, '{'{-25'd378164}}, '{'{25'd2100913}}, '{'{25'd2016876}}, '{'{-25'd588256}}, '{'{-25'd336146}}, '{'{-25'd756329}}, '{'{25'd2058894}}, '{'{25'd1806785}}, '{'{-25'd840365}}, '{'{25'd2353022}}, '{'{-25'd3949716}}, '{'{25'd1890821}}, '{'{-25'd1092475}}, '{'{-25'd756329}}, '{'{-25'd1344584}}, '{'{-25'd840365}}, '{'{-25'd5336318}}, '{'{25'd1512657}}, '{'{25'd1344584}}, '{'{-25'd1344584}}, '{'{25'd2479077}}},
    '{'{'{25'd2023241}}, '{'{-25'd1416268}}, '{'{25'd303486}}, '{'{-25'd3490090}}, '{'{-25'd556391}}, '{'{-25'd4097062}}, '{'{-25'd2478470}}, '{'{25'd1669173}}, '{'{-25'd2124403}}, '{'{-25'd1213944}}, '{'{-25'd1011620}}, '{'{25'd252905}}, '{'{-25'd4046481}}, '{'{-25'd2832537}}, '{'{-25'd1820917}}, '{'{-25'd2883118}}, '{'{-25'd6474370}}, '{'{25'd303486}}, '{'{25'd0}}, '{'{25'd0}}, '{'{25'd505810}}, '{'{25'd5108682}}, '{'{-25'd404648}}, '{'{25'd5867398}}, '{'{-25'd101162}}, '{'{-25'd2073822}}, '{'{25'd1922079}}, '{'{25'd5311007}}, '{'{25'd5462750}}, '{'{-25'd50581}}, '{'{-25'd606972}}, '{'{-25'd1618592}}, '{'{25'd2174984}}, '{'{-25'd1517430}}, '{'{-25'd3490090}}, '{'{-25'd2023241}}, '{'{-25'd3136023}}, '{'{-25'd961039}}, '{'{25'd1315106}}, '{'{-25'd1112782}}, '{'{25'd354067}}, '{'{25'd1669173}}, '{'{25'd1922079}}, '{'{25'd758715}}, '{'{-25'd1922079}}, '{'{25'd1011620}}, '{'{-25'd1062201}}, '{'{25'd1011620}}, '{'{-25'd2427889}}, '{'{-25'd455229}}, '{'{25'd1770336}}, '{'{-25'd1112782}}, '{'{25'd910458}}, '{'{25'd505810}}, '{'{-25'd1568011}}, '{'{25'd1466849}}, '{'{-25'd809296}}, '{'{25'd1972660}}, '{'{25'd404648}}, '{'{25'd5563912}}, '{'{-25'd1112782}}, '{'{25'd2276146}}, '{'{-25'd1011620}}, '{'{25'd1517430}}},
    '{'{'{-25'd2473133}}, '{'{25'd1723699}}, '{'{25'd2585548}}, '{'{-25'd2173359}}, '{'{25'd674491}}, '{'{25'd1873586}}, '{'{25'd3072680}}, '{'{-25'd1199095}}, '{'{25'd1086680}}, '{'{-25'd1274038}}, '{'{-25'd374717}}, '{'{25'd37472}}, '{'{-25'd1161623}}, '{'{25'd412189}}, '{'{25'd449661}}, '{'{-25'd2210831}}, '{'{-25'd1648755}}, '{'{-25'd1386453}}, '{'{-25'd1536340}}, '{'{25'd2210831}}, '{'{-25'd74943}}, '{'{-25'd149887}}, '{'{-25'd2098416}}, '{'{-25'd1798642}}, '{'{-25'd2435661}}, '{'{-25'd149887}}, '{'{25'd1986001}}, '{'{25'd1536340}}, '{'{25'd4758907}}, '{'{25'd224830}}, '{'{25'd74943}}, '{'{25'd412189}}, '{'{25'd487132}}, '{'{25'd1536340}}, '{'{-25'd1274038}}, '{'{25'd2173359}}, '{'{-25'd786906}}, '{'{25'd74943}}, '{'{-25'd74943}}, '{'{25'd2098416}}, '{'{-25'd1573812}}, '{'{25'd2510605}}, '{'{25'd2173359}}, '{'{25'd0}}, '{'{-25'd711962}}, '{'{-25'd1498868}}, '{'{25'd899321}}, '{'{25'd2360718}}, '{'{-25'd2660491}}, '{'{25'd1536340}}, '{'{-25'd337245}}, '{'{25'd1011736}}, '{'{25'd1611284}}, '{'{25'd2173359}}, '{'{-25'd1573812}}, '{'{25'd1461397}}, '{'{25'd112415}}, '{'{-25'd936793}}, '{'{-25'd149887}}, '{'{25'd4121888}}, '{'{25'd1423925}}, '{'{25'd2323246}}, '{'{25'd674491}}, '{'{-25'd2135887}}},
    '{'{'{25'd799427}}, '{'{25'd1065902}}, '{'{25'd799427}}, '{'{25'd2339063}}, '{'{-25'd177650}}, '{'{-25'd799427}}, '{'{25'd473734}}, '{'{25'd384909}}, '{'{25'd710601}}, '{'{-25'd858643}}, '{'{25'd2102196}}, '{'{25'd1806112}}, '{'{-25'd59217}}, '{'{-25'd2339063}}, '{'{25'd177650}}, '{'{25'd148042}}, '{'{25'd473734}}, '{'{-25'd621776}}, '{'{-25'd2931231}}, '{'{25'd236867}}, '{'{25'd740210}}, '{'{25'd1894937}}, '{'{-25'd1510028}}, '{'{-25'd1095511}}, '{'{25'd148042}}, '{'{-25'd2013371}}, '{'{-25'd829035}}, '{'{-25'd621776}}, '{'{-25'd355301}}, '{'{25'd2427888}}, '{'{25'd266476}}, '{'{-25'd1598853}}, '{'{25'd118434}}, '{'{-25'd947469}}, '{'{25'd977077}}, '{'{25'd2250238}}, '{'{25'd2309455}}, '{'{-25'd740210}}, '{'{25'd1065902}}, '{'{25'd2279846}}, '{'{25'd1243553}}, '{'{-25'd1332378}}, '{'{-25'd858643}}, '{'{25'd1480420}}, '{'{-25'd2131804}}, '{'{-25'd88825}}, '{'{25'd384909}}, '{'{25'd1687679}}, '{'{25'd3375357}}, '{'{25'd621776}}, '{'{25'd1243553}}, '{'{25'd1835721}}, '{'{-25'd1006685}}, '{'{-25'd3168098}}, '{'{-25'd3760266}}, '{'{25'd1717287}}, '{'{25'd1243553}}, '{'{25'd148042}}, '{'{25'd2516714}}, '{'{-25'd2427888}}, '{'{25'd977077}}, '{'{25'd1539637}}, '{'{25'd2723972}}, '{'{-25'd1658070}}},
    '{'{'{-25'd1743522}}, '{'{25'd2122548}}, '{'{25'd4472512}}, '{'{25'd1819327}}, '{'{-25'd720150}}, '{'{-25'd947566}}, '{'{-25'd379026}}, '{'{-25'd1212885}}, '{'{-25'd1099177}}, '{'{-25'd644345}}, '{'{-25'd1743522}}, '{'{-25'd644345}}, '{'{-25'd720150}}, '{'{25'd2160451}}, '{'{25'd909664}}, '{'{25'd1250787}}, '{'{-25'd2046743}}, '{'{25'd947566}}, '{'{25'd758053}}, '{'{-25'd2160451}}, '{'{25'd1061274}}, '{'{25'd1250787}}, '{'{-25'd682248}}, '{'{-25'd1591911}}, '{'{-25'd2274159}}, '{'{25'd530637}}, '{'{-25'd2312062}}, '{'{25'd1667717}}, '{'{-25'd189513}}, '{'{25'd2084646}}, '{'{-25'd1516106}}, '{'{25'd720150}}, '{'{25'd492734}}, '{'{-25'd682248}}, '{'{-25'd1819327}}, '{'{25'd2160451}}, '{'{-25'd1933035}}, '{'{25'd1629814}}, '{'{25'd720150}}, '{'{-25'd1895132}}, '{'{25'd2653185}}, '{'{-25'd3449141}}, '{'{-25'd151611}}, '{'{25'd1667717}}, '{'{-25'd37903}}, '{'{25'd1478203}}, '{'{25'd2349964}}, '{'{25'd1516106}}, '{'{25'd4813636}}, '{'{-25'd227416}}, '{'{25'd833858}}, '{'{25'd947566}}, '{'{25'd1288690}}, '{'{25'd2766893}}, '{'{-25'd189513}}, '{'{-25'd1326593}}, '{'{25'd492734}}, '{'{25'd1364495}}, '{'{-25'd2160451}}, '{'{25'd1478203}}, '{'{-25'd795956}}, '{'{-25'd530637}}, '{'{25'd2463672}}, '{'{-25'd1667717}}},
    '{'{'{-25'd2264554}}, '{'{25'd226455}}, '{'{-25'd543493}}, '{'{25'd1494606}}, '{'{-25'd1449314}}, '{'{25'd1902225}}, '{'{25'd3170375}}, '{'{25'd226455}}, '{'{-25'd860530}}, '{'{25'd498202}}, '{'{-25'd2128681}}, '{'{25'd1811643}}, '{'{-25'd1992807}}, '{'{-25'd860530}}, '{'{25'd1766352}}, '{'{25'd2626882}}, '{'{-25'd1132277}}, '{'{25'd226455}}, '{'{-25'd1766352}}, '{'{25'd498202}}, '{'{25'd90582}}, '{'{25'd3306249}}, '{'{25'd679366}}, '{'{25'd905822}}, '{'{25'd2309845}}, '{'{25'd2400427}}, '{'{-25'd951113}}, '{'{25'd2219263}}, '{'{25'd4936727}}, '{'{25'd1992807}}, '{'{25'd407620}}, '{'{25'd1132277}}, '{'{25'd860530}}, '{'{25'd498202}}, '{'{-25'd1222859}}, '{'{-25'd634075}}, '{'{-25'd2898629}}, '{'{25'd634075}}, '{'{25'd1630479}}, '{'{-25'd1222859}}, '{'{25'd498202}}, '{'{25'd860530}}, '{'{-25'd1358732}}, '{'{-25'd1766352}}, '{'{25'd2219263}}, '{'{25'd1449314}}, '{'{-25'd452911}}, '{'{25'd2173972}}, '{'{25'd5751967}}, '{'{-25'd2038098}}, '{'{25'd2038098}}, '{'{25'd951113}}, '{'{-25'd1539897}}, '{'{25'd1902225}}, '{'{-25'd3623286}}, '{'{-25'd1494606}}, '{'{-25'd1449314}}, '{'{25'd1449314}}, '{'{-25'd1675770}}, '{'{-25'd2762756}}, '{'{-25'd1856934}}, '{'{25'd1494606}}, '{'{25'd1449314}}, '{'{25'd2038098}}},
    '{'{'{-25'd1294189}}, '{'{25'd1119298}}, '{'{-25'd174890}}, '{'{25'd1678947}}, '{'{-25'd979386}}, '{'{25'd2238597}}, '{'{25'd1049342}}, '{'{-25'd1504057}}, '{'{-25'd1014364}}, '{'{25'd2098684}}, '{'{25'd419737}}, '{'{25'd0}}, '{'{-25'd1259211}}, '{'{25'd1853838}}, '{'{-25'd69956}}, '{'{-25'd1539035}}, '{'{25'd1189254}}, '{'{-25'd1469079}}, '{'{25'd3287939}}, '{'{-25'd839474}}, '{'{-25'd1853838}}, '{'{-25'd4477193}}, '{'{-25'd2308553}}, '{'{-25'd524671}}, '{'{25'd2903180}}, '{'{25'd2238597}}, '{'{-25'd1958772}}, '{'{25'd4232347}}, '{'{25'd3113048}}, '{'{-25'd1329167}}, '{'{-25'd1434101}}, '{'{-25'd1958772}}, '{'{-25'd1608991}}, '{'{25'd1748904}}, '{'{-25'd2063706}}, '{'{25'd1853838}}, '{'{-25'd454715}}, '{'{-25'd594627}}, '{'{-25'd209868}}, '{'{-25'd979386}}, '{'{-25'd1154276}}, '{'{25'd0}}, '{'{-25'd559649}}, '{'{25'd1329167}}, '{'{25'd1678947}}, '{'{-25'd279825}}, '{'{-25'd559649}}, '{'{25'd804496}}, '{'{-25'd1364145}}, '{'{-25'd1364145}}, '{'{25'd594627}}, '{'{25'd279825}}, '{'{-25'd454715}}, '{'{-25'd3602741}}, '{'{-25'd3008114}}, '{'{-25'd1713925}}, '{'{25'd1329167}}, '{'{-25'd2343531}}, '{'{25'd2063706}}, '{'{-25'd1574013}}, '{'{-25'd454715}}, '{'{25'd1084320}}, '{'{25'd279825}}, '{'{-25'd1364145}}},
    '{'{'{-25'd69280}}, '{'{25'd1177757}}, '{'{25'd207839}}, '{'{-25'd1801276}}, '{'{25'd2632634}}, '{'{25'd2424794}}, '{'{-25'd969918}}, '{'{25'd1454876}}, '{'{25'd762078}}, '{'{-25'd1247037}}, '{'{25'd1454876}}, '{'{-25'd1108477}}, '{'{25'd415679}}, '{'{25'd2632634}}, '{'{25'd1385597}}, '{'{-25'd8867818}}, '{'{25'd138560}}, '{'{-25'd1247037}}, '{'{25'd1316317}}, '{'{-25'd1731996}}, '{'{25'd2147675}}, '{'{-25'd415679}}, '{'{25'd554239}}, '{'{25'd3741111}}, '{'{25'd1039197}}, '{'{25'd1316317}}, '{'{25'd1247037}}, '{'{25'd4087510}}, '{'{25'd1731996}}, '{'{25'd138560}}, '{'{25'd1801276}}, '{'{25'd2078395}}, '{'{-25'd1108477}}, '{'{25'd415679}}, '{'{25'd3186872}}, '{'{25'd207839}}, '{'{25'd277119}}, '{'{-25'd277119}}, '{'{-25'd1662716}}, '{'{25'd138560}}, '{'{25'd4572469}}, '{'{25'd2355514}}, '{'{-25'd346399}}, '{'{25'd1247037}}, '{'{-25'd1939835}}, '{'{25'd277119}}, '{'{-25'd692798}}, '{'{25'd2424794}}, '{'{-25'd3533271}}, '{'{-25'd969918}}, '{'{25'd2009115}}, '{'{-25'd2078395}}, '{'{-25'd2009115}}, '{'{25'd6581584}}, '{'{25'd2286234}}, '{'{25'd1177757}}, '{'{-25'd2147675}}, '{'{-25'd2286234}}, '{'{25'd1939835}}, '{'{25'd4226070}}, '{'{25'd2286234}}, '{'{25'd1316317}}, '{'{25'd3741111}}, '{'{-25'd1939835}}},
    '{'{'{25'd2263812}}, '{'{25'd1890400}}, '{'{25'd1073561}}, '{'{25'd1727032}}, '{'{25'd1493649}}, '{'{25'd23338}}, '{'{25'd2567210}}, '{'{25'd1493649}}, '{'{-25'd1283605}}, '{'{25'd2263812}}, '{'{25'd1750370}}, '{'{25'd350074}}, '{'{-25'd840178}}, '{'{-25'd466765}}, '{'{-25'd2217136}}, '{'{-25'd46677}}, '{'{-25'd116691}}, '{'{-25'd1937077}}, '{'{25'd933531}}, '{'{25'd1423635}}, '{'{25'd1050222}}, '{'{25'd1120237}}, '{'{25'd1867062}}, '{'{-25'd700148}}, '{'{25'd256721}}, '{'{25'd186706}}, '{'{25'd2333827}}, '{'{-25'd466765}}, '{'{-25'd2193798}}, '{'{25'd490104}}, '{'{25'd1003546}}, '{'{25'd1516988}}, '{'{-25'd1213590}}, '{'{-25'd1680356}}, '{'{-25'd1283605}}, '{'{25'd490104}}, '{'{-25'd1797047}}, '{'{25'd1890400}}, '{'{-25'd1493649}}, '{'{25'd2217136}}, '{'{25'd46677}}, '{'{-25'd723486}}, '{'{25'd1283605}}, '{'{25'd1913738}}, '{'{-25'd1937077}}, '{'{-25'd583457}}, '{'{25'd700148}}, '{'{25'd2147121}}, '{'{25'd1587003}}, '{'{-25'd1890400}}, '{'{25'd303398}}, '{'{25'd303398}}, '{'{-25'd2380504}}, '{'{-25'd2543872}}, '{'{-25'd303398}}, '{'{25'd1376958}}, '{'{25'd816840}}, '{'{-25'd2193798}}, '{'{25'd1773709}}, '{'{25'd583457}}, '{'{-25'd1470311}}, '{'{-25'd443427}}, '{'{25'd2963961}}, '{'{25'd326736}}},
    '{'{'{25'd314179}}, '{'{25'd1832713}}, '{'{25'd2565799}}, '{'{-25'd837812}}, '{'{-25'd3089431}}, '{'{25'd1466171}}, '{'{25'd1256718}}, '{'{-25'd1151991}}, '{'{25'd785449}}, '{'{-25'd2042166}}, '{'{-25'd2408709}}, '{'{-25'd1832713}}, '{'{-25'd366543}}, '{'{25'd1989803}}, '{'{-25'd314179}}, '{'{25'd2094529}}, '{'{-25'd1989803}}, '{'{-25'd575996}}, '{'{-25'd1727987}}, '{'{25'd314179}}, '{'{-25'd2094529}}, '{'{-25'd1780350}}, '{'{-25'd1727987}}, '{'{25'd6650131}}, '{'{25'd157090}}, '{'{-25'd2042166}}, '{'{-25'd2146893}}, '{'{25'd3665427}}, '{'{25'd1047265}}, '{'{25'd1623260}}, '{'{-25'd1518534}}, '{'{25'd2303982}}, '{'{25'd1727987}}, '{'{-25'd1570897}}, '{'{-25'd52363}}, '{'{-25'd314179}}, '{'{-25'd1675624}}, '{'{25'd1675624}}, '{'{25'd628359}}, '{'{25'd1309081}}, '{'{25'd2879978}}, '{'{-25'd1780350}}, '{'{25'd2356346}}, '{'{-25'd942538}}, '{'{25'd2094529}}, '{'{-25'd1832713}}, '{'{25'd471269}}, '{'{25'd3770153}}, '{'{25'd366543}}, '{'{25'd837812}}, '{'{-25'd733085}}, '{'{-25'd1989803}}, '{'{25'd2827615}}, '{'{-25'd1780350}}, '{'{-25'd680722}}, '{'{-25'd1256718}}, '{'{25'd1518534}}, '{'{-25'd314179}}, '{'{-25'd314179}}, '{'{25'd5288687}}, '{'{25'd1309081}}, '{'{-25'd4241422}}, '{'{-25'd1256718}}, '{'{25'd1309081}}},
    '{'{'{25'd1049551}}, '{'{-25'd185215}}, '{'{-25'd926075}}, '{'{-25'd802598}}, '{'{25'd493906}}, '{'{25'd555645}}, '{'{25'd864336}}, '{'{25'd1234766}}, '{'{25'd1852149}}, '{'{25'd1543458}}, '{'{25'd1543458}}, '{'{25'd555645}}, '{'{-25'd4445158}}, '{'{25'd2839962}}, '{'{-25'd1852149}}, '{'{25'd1358243}}, '{'{25'd987813}}, '{'{25'd432168}}, '{'{25'd1852149}}, '{'{-25'd926075}}, '{'{-25'd679121}}, '{'{-25'd2222579}}, '{'{-25'd617383}}, '{'{-25'd987813}}, '{'{-25'd1481719}}, '{'{-25'd1975626}}, '{'{25'd1790411}}, '{'{25'd2284317}}, '{'{25'd493906}}, '{'{-25'd1543458}}, '{'{-25'd802598}}, '{'{-25'd1728673}}, '{'{25'd555645}}, '{'{-25'd2037364}}, '{'{25'd2037364}}, '{'{25'd308692}}, '{'{-25'd1358243}}, '{'{25'd2407794}}, '{'{-25'd1605196}}, '{'{25'd926075}}, '{'{-25'd987813}}, '{'{-25'd1481719}}, '{'{25'd1049551}}, '{'{-25'd308692}}, '{'{-25'd1173028}}, '{'{25'd1358243}}, '{'{-25'd1358243}}, '{'{25'd1296504}}, '{'{-25'd2593009}}, '{'{-25'd432168}}, '{'{25'd2346056}}, '{'{25'd185215}}, '{'{-25'd370430}}, '{'{-25'd61738}}, '{'{25'd5494709}}, '{'{25'd1296504}}, '{'{-25'd2407794}}, '{'{25'd1543458}}, '{'{-25'd617383}}, '{'{-25'd7902503}}, '{'{25'd2160841}}, '{'{-25'd1358243}}, '{'{-25'd1605196}}, '{'{-25'd1975626}}},
    '{'{'{25'd0}}, '{'{-25'd990850}}, '{'{25'd1378574}}, '{'{25'd1723218}}, '{'{25'd172322}}, '{'{-25'd2627907}}, '{'{-25'd1766298}}, '{'{25'd215402}}, '{'{-25'd2154022}}, '{'{-25'd1033931}}, '{'{25'd1335494}}, '{'{-25'd258483}}, '{'{-25'd430804}}, '{'{-25'd129241}}, '{'{-25'd516965}}, '{'{-25'd603126}}, '{'{25'd947770}}, '{'{-25'd1852459}}, '{'{25'd818528}}, '{'{-25'd775448}}, '{'{-25'd689287}}, '{'{-25'd560046}}, '{'{25'd861609}}, '{'{25'd5471216}}, '{'{-25'd1249333}}, '{'{25'd2369424}}, '{'{25'd1033931}}, '{'{25'd4825009}}, '{'{25'd2541746}}, '{'{25'd86161}}, '{'{-25'd516965}}, '{'{-25'd732367}}, '{'{-25'd430804}}, '{'{-25'd689287}}, '{'{25'd4480366}}, '{'{-25'd473885}}, '{'{-25'd1163172}}, '{'{25'd2843309}}, '{'{-25'd1378574}}, '{'{25'd1378574}}, '{'{25'd172322}}, '{'{25'd2369424}}, '{'{-25'd301563}}, '{'{25'd1421655}}, '{'{25'd43080}}, '{'{-25'd732367}}, '{'{25'd560046}}, '{'{25'd1292413}}, '{'{25'd1809379}}, '{'{25'd1077011}}, '{'{-25'd1507815}}, '{'{-25'd516965}}, '{'{25'd1335494}}, '{'{-25'd5212733}}, '{'{25'd258483}}, '{'{25'd2326344}}, '{'{-25'd2067861}}, '{'{25'd2067861}}, '{'{25'd43080}}, '{'{25'd1680137}}, '{'{25'd43080}}, '{'{-25'd1593976}}, '{'{25'd1507815}}, '{'{25'd2541746}}},
    '{'{'{-25'd2177208}}, '{'{25'd2305279}}, '{'{25'd3778095}}, '{'{25'd1792994}}, '{'{25'd2017119}}, '{'{-25'd672373}}, '{'{25'd1408781}}, '{'{25'd1889048}}, '{'{-25'd1152639}}, '{'{-25'd1440799}}, '{'{25'd352195}}, '{'{25'd1248693}}, '{'{-25'd3618007}}, '{'{-25'd192107}}, '{'{25'd128071}}, '{'{-25'd736408}}, '{'{-25'd2241243}}, '{'{25'd128071}}, '{'{-25'd4098273}}, '{'{-25'd1632906}}, '{'{-25'd32018}}, '{'{-25'd1472817}}, '{'{-25'd2049137}}, '{'{-25'd768426}}, '{'{-25'd1664923}}, '{'{-25'd1504835}}, '{'{-25'd2145190}}, '{'{25'd608337}}, '{'{-25'd704391}}, '{'{-25'd1248693}}, '{'{25'd2209225}}, '{'{25'd2049137}}, '{'{-25'd1344746}}, '{'{-25'd1504835}}, '{'{25'd192107}}, '{'{25'd1184657}}, '{'{25'd1312728}}, '{'{25'd288160}}, '{'{-25'd2017119}}, '{'{-25'd2081154}}, '{'{-25'd992551}}, '{'{25'd1536852}}, '{'{-25'd1152639}}, '{'{25'd768426}}, '{'{25'd2305279}}, '{'{25'd224124}}, '{'{-25'd960533}}, '{'{-25'd1088604}}, '{'{-25'd480266}}, '{'{25'd544302}}, '{'{25'd768426}}, '{'{-25'd1728959}}, '{'{-25'd1857030}}, '{'{25'd3618007}}, '{'{25'd0}}, '{'{25'd2561421}}, '{'{25'd1056586}}, '{'{25'd2049137}}, '{'{25'd1600888}}, '{'{-25'd640355}}, '{'{25'd128071}}, '{'{-25'd1664923}}, '{'{-25'd736408}}, '{'{-25'd1953083}}},
    '{'{'{25'd164103}}, '{'{-25'd1936416}}, '{'{-25'd1115901}}, '{'{-25'd2133340}}, '{'{-25'd1411286}}, '{'{-25'd98462}}, '{'{25'd3314882}}, '{'{25'd623592}}, '{'{25'd1641031}}, '{'{-25'd32821}}, '{'{-25'd295386}}, '{'{-25'd1050260}}, '{'{-25'd2494367}}, '{'{-25'd2363084}}, '{'{-25'd557950}}, '{'{-25'd361027}}, '{'{25'd2100519}}, '{'{25'd2166160}}, '{'{-25'd65641}}, '{'{25'd2133340}}, '{'{25'd1837954}}, '{'{25'd689233}}, '{'{-25'd1608210}}, '{'{-25'd3905653}}, '{'{25'd656412}}, '{'{25'd1575389}}, '{'{-25'd65641}}, '{'{-25'd4102577}}, '{'{25'd131282}}, '{'{-25'd951798}}, '{'{25'd2592828}}, '{'{25'd2330264}}, '{'{25'd0}}, '{'{-25'd2297443}}, '{'{-25'd1247183}}, '{'{-25'd853336}}, '{'{25'd1181542}}, '{'{25'd2330264}}, '{'{25'd1378466}}, '{'{25'd1411286}}, '{'{-25'd2461546}}, '{'{25'd2264622}}, '{'{-25'd98462}}, '{'{25'd1214363}}, '{'{-25'd1312825}}, '{'{25'd2363084}}, '{'{25'd1805134}}, '{'{-25'd1378466}}, '{'{-25'd2986676}}, '{'{25'd754874}}, '{'{-25'd32821}}, '{'{25'd1181542}}, '{'{25'd2067699}}, '{'{25'd4168218}}, '{'{-25'd3840012}}, '{'{-25'd1083080}}, '{'{25'd1870775}}, '{'{25'd2297443}}, '{'{-25'd131282}}, '{'{-25'd1345645}}, '{'{25'd2625649}}, '{'{-25'd2166160}}, '{'{-25'd3249241}}, '{'{-25'd525130}}},
    '{'{'{-25'd293963}}, '{'{-25'd1665788}}, '{'{-25'd1665788}}, '{'{-25'd391950}}, '{'{25'd293963}}, '{'{25'd1796438}}, '{'{25'd457275}}, '{'{-25'd1992413}}, '{'{25'd391950}}, '{'{25'd1633125}}, '{'{25'd1077863}}, '{'{25'd2482351}}, '{'{-25'd1045200}}, '{'{-25'd4180801}}, '{'{-25'd1208513}}, '{'{25'd718575}}, '{'{-25'd1894426}}, '{'{-25'd2482351}}, '{'{25'd522600}}, '{'{25'd293963}}, '{'{25'd816563}}, '{'{25'd2090401}}, '{'{-25'd1698450}}, '{'{-25'd1306500}}, '{'{-25'd2319038}}, '{'{-25'd1273838}}, '{'{25'd2221051}}, '{'{25'd1763776}}, '{'{-25'd2351701}}, '{'{25'd2808976}}, '{'{-25'd1698450}}, '{'{-25'd2025076}}, '{'{25'd32663}}, '{'{-25'd555263}}, '{'{25'd2351701}}, '{'{-25'd1796438}}, '{'{-25'd1502475}}, '{'{25'd130650}}, '{'{25'd130650}}, '{'{25'd555263}}, '{'{25'd2123063}}, '{'{-25'd1175850}}, '{'{25'd979875}}, '{'{-25'd1992413}}, '{'{25'd424613}}, '{'{25'd2808976}}, '{'{-25'd1796438}}, '{'{25'd2090401}}, '{'{-25'd1535138}}, '{'{-25'd489938}}, '{'{-25'd228638}}, '{'{-25'd685913}}, '{'{-25'd620588}}, '{'{25'd1763776}}, '{'{25'd1175850}}, '{'{-25'd2645663}}, '{'{-25'd1861763}}, '{'{-25'd1763776}}, '{'{-25'd65325}}, '{'{-25'd1371825}}, '{'{-25'd2417026}}, '{'{25'd2678326}}, '{'{-25'd2319038}}, '{'{25'd979875}}},
    '{'{'{-25'd2190215}}, '{'{-25'd2570150}}, '{'{25'd1519741}}, '{'{25'd1407995}}, '{'{25'd692823}}, '{'{-25'd1296250}}, '{'{-25'd1452694}}, '{'{25'd1989073}}, '{'{-25'd759871}}, '{'{25'd2123168}}, '{'{25'd223491}}, '{'{-25'd1095108}}, '{'{-25'd178793}}, '{'{25'd290539}}, '{'{25'd1072758}}, '{'{-25'd1854978}}, '{'{25'd1072758}}, '{'{25'd1363297}}, '{'{-25'd201142}}, '{'{25'd134095}}, '{'{25'd2838340}}, '{'{-25'd1609138}}, '{'{25'd1787931}}, '{'{-25'd469332}}, '{'{25'd1989073}}, '{'{25'd1854978}}, '{'{25'd2346659}}, '{'{25'd737521}}, '{'{25'd961013}}, '{'{25'd581077}}, '{'{-25'd1743232}}, '{'{-25'd1899676}}, '{'{-25'd2100819}}, '{'{25'd1542090}}, '{'{25'd916315}}, '{'{-25'd1653836}}, '{'{25'd1989073}}, '{'{25'd2547801}}, '{'{-25'd1095108}}, '{'{-25'd1877327}}, '{'{25'd1430345}}, '{'{-25'd871616}}, '{'{-25'd2324310}}, '{'{25'd335237}}, '{'{-25'd2458405}}, '{'{-25'd648125}}, '{'{25'd223491}}, '{'{-25'd2793642}}, '{'{25'd1340948}}, '{'{-25'd1273901}}, '{'{-25'd2681896}}, '{'{25'd2011422}}, '{'{25'd1899676}}, '{'{25'd2838340}}, '{'{25'd826918}}, '{'{-25'd849267}}, '{'{25'd2324310}}, '{'{25'd1787931}}, '{'{-25'd2056120}}, '{'{25'd2033771}}, '{'{-25'd1698534}}, '{'{25'd156444}}, '{'{-25'd1854978}}, '{'{-25'd1050409}}},
    '{'{'{-25'd1717606}}, '{'{25'd1679437}}, '{'{25'd3511550}}, '{'{-25'd1488592}}, '{'{-25'd114507}}, '{'{-25'd381690}}, '{'{-25'd381690}}, '{'{25'd2175635}}, '{'{25'd2290142}}, '{'{-25'd38169}}, '{'{-25'd877888}}, '{'{-25'd1068733}}, '{'{-25'd2137465}}, '{'{-25'd1755775}}, '{'{25'd1335916}}, '{'{25'd916057}}, '{'{25'd2519156}}, '{'{-25'd801550}}, '{'{-25'd1564930}}, '{'{25'd190845}}, '{'{-25'd2328311}}, '{'{25'd152676}}, '{'{25'd76338}}, '{'{25'd877888}}, '{'{-25'd38169}}, '{'{-25'd190845}}, '{'{-25'd648873}}, '{'{-25'd725212}}, '{'{25'd458028}}, '{'{25'd1259578}}, '{'{25'd839719}}, '{'{-25'd839719}}, '{'{25'd2595494}}, '{'{-25'd1221409}}, '{'{25'd2137465}}, '{'{25'd1068733}}, '{'{25'd1908451}}, '{'{25'd1030564}}, '{'{25'd2519156}}, '{'{25'd419859}}, '{'{25'd1450423}}, '{'{-25'd1755775}}, '{'{-25'd2251973}}, '{'{-25'd114507}}, '{'{25'd1717606}}, '{'{-25'd916057}}, '{'{-25'd2939015}}, '{'{-25'd1335916}}, '{'{-25'd2595494}}, '{'{25'd1870282}}, '{'{25'd2366480}}, '{'{25'd305352}}, '{'{-25'd2290142}}, '{'{25'd0}}, '{'{-25'd4847466}}, '{'{25'd343521}}, '{'{-25'd763381}}, '{'{25'd229014}}, '{'{25'd305352}}, '{'{25'd1870282}}, '{'{-25'd305352}}, '{'{25'd2137465}}, '{'{25'd3778734}}, '{'{-25'd877888}}},
    '{'{'{25'd1376320}}, '{'{25'd2395817}}, '{'{25'd1733144}}, '{'{25'd1631195}}, '{'{-25'd866572}}, '{'{25'd1988018}}, '{'{-25'd1376320}}, '{'{25'd1937044}}, '{'{25'd1784119}}, '{'{-25'd2140943}}, '{'{25'd815597}}, '{'{25'd1733144}}, '{'{-25'd1631195}}, '{'{-25'd866572}}, '{'{25'd1223396}}, '{'{25'd6473804}}, '{'{25'd713648}}, '{'{25'd1376320}}, '{'{-25'd1886069}}, '{'{25'd1937044}}, '{'{-25'd356824}}, '{'{-25'd2242893}}, '{'{25'd2140943}}, '{'{-25'd713648}}, '{'{-25'd50975}}, '{'{-25'd866572}}, '{'{-25'd2395817}}, '{'{-25'd1529245}}, '{'{25'd611698}}, '{'{25'd1886069}}, '{'{-25'd2344842}}, '{'{25'd1733144}}, '{'{-25'd1070471}}, '{'{-25'd917547}}, '{'{-25'd407799}}, '{'{25'd101950}}, '{'{25'd713648}}, '{'{-25'd407799}}, '{'{25'd662673}}, '{'{25'd1886069}}, '{'{25'd2242893}}, '{'{25'd1478270}}, '{'{25'd1427295}}, '{'{-25'd1019497}}, '{'{-25'd1223396}}, '{'{-25'd611698}}, '{'{-25'd1274371}}, '{'{-25'd407799}}, '{'{25'd1937044}}, '{'{25'd407799}}, '{'{25'd764622}}, '{'{25'd254874}}, '{'{-25'd1376320}}, '{'{25'd407799}}, '{'{-25'd2242893}}, '{'{-25'd764622}}, '{'{25'd917547}}, '{'{-25'd2344842}}, '{'{25'd1325346}}, '{'{-25'd4995534}}, '{'{-25'd2293867}}, '{'{25'd1682169}}, '{'{25'd815597}}, '{'{25'd1988018}}},
    '{'{'{-25'd1372685}}, '{'{-25'd492759}}, '{'{25'd1126305}}, '{'{25'd844729}}, '{'{25'd774335}}, '{'{-25'd703941}}, '{'{25'd3238128}}, '{'{25'd774335}}, '{'{-25'd703941}}, '{'{25'd0}}, '{'{-25'd1795049}}, '{'{-25'd1020714}}, '{'{25'd70394}}, '{'{25'd1865443}}, '{'{25'd175985}}, '{'{25'd739138}}, '{'{-25'd985517}}, '{'{25'd809532}}, '{'{25'd1478276}}, '{'{25'd1055911}}, '{'{25'd1971035}}, '{'{-25'd387167}}, '{'{-25'd2006232}}, '{'{25'd492759}}, '{'{-25'd527956}}, '{'{-25'd1900640}}, '{'{-25'd1020714}}, '{'{-25'd1724655}}, '{'{25'd4470025}}, '{'{-25'd598350}}, '{'{-25'd1161502}}, '{'{-25'd527956}}, '{'{25'd1548670}}, '{'{25'd1267094}}, '{'{25'd1267094}}, '{'{25'd70394}}, '{'{25'd1020714}}, '{'{-25'd2182217}}, '{'{25'd1055911}}, '{'{-25'd1055911}}, '{'{-25'd316773}}, '{'{-25'd35197}}, '{'{25'd1759852}}, '{'{25'd2076626}}, '{'{25'd1865443}}, '{'{25'd1372685}}, '{'{-25'd2076626}}, '{'{-25'd1619064}}, '{'{-25'd1689458}}, '{'{25'd1478276}}, '{'{25'd739138}}, '{'{25'd563153}}, '{'{25'd2006232}}, '{'{-25'd2815764}}, '{'{25'd2393399}}, '{'{25'd2006232}}, '{'{-25'd2076626}}, '{'{25'd915123}}, '{'{-25'd1126305}}, '{'{25'd3519704}}, '{'{25'd0}}, '{'{25'd246379}}, '{'{-25'd703941}}, '{'{25'd1724655}}},
    '{'{'{25'd1131330}}, '{'{-25'd1759847}}, '{'{25'd911349}}, '{'{-25'd1351311}}, '{'{-25'd1037053}}, '{'{25'd2325512}}, '{'{25'd3991082}}, '{'{25'd502813}}, '{'{-25'd439962}}, '{'{-25'd2042680}}, '{'{-25'd2042680}}, '{'{-25'd1351311}}, '{'{-25'd2859751}}, '{'{-25'd2482641}}, '{'{25'd1319885}}, '{'{-25'd1822699}}, '{'{25'd659943}}, '{'{25'd2231235}}, '{'{25'd942775}}, '{'{25'd2042680}}, '{'{25'd2451215}}, '{'{25'd1854124}}, '{'{25'd125703}}, '{'{25'd408536}}, '{'{25'd62852}}, '{'{25'd722794}}, '{'{25'd1225608}}, '{'{-25'd628517}}, '{'{25'd62852}}, '{'{-25'd691368}}, '{'{25'd2356938}}, '{'{25'd1445589}}, '{'{25'd251407}}, '{'{25'd1508440}}, '{'{25'd1319885}}, '{'{25'd251407}}, '{'{-25'd2074105}}, '{'{25'd2262660}}, '{'{-25'd1131330}}, '{'{-25'd1634144}}, '{'{25'd1037053}}, '{'{25'd2482641}}, '{'{-25'd1979828}}, '{'{-25'd2074105}}, '{'{-25'd848498}}, '{'{25'd2199809}}, '{'{25'd502813}}, '{'{-25'd219981}}, '{'{-25'd188555}}, '{'{25'd1539866}}, '{'{25'd722794}}, '{'{25'd377110}}, '{'{-25'd1634144}}, '{'{25'd2042680}}, '{'{-25'd1351311}}, '{'{-25'd1539866}}, '{'{25'd2168383}}, '{'{-25'd1508440}}, '{'{25'd2042680}}, '{'{25'd848498}}, '{'{-25'd1822699}}, '{'{25'd1005627}}, '{'{-25'd1728421}}, '{'{-25'd125703}}},
    '{'{'{25'd1760733}}, '{'{-25'd1844577}}, '{'{-25'd922289}}, '{'{-25'd1383433}}, '{'{-25'd1467277}}, '{'{-25'd2012266}}, '{'{-25'd754600}}, '{'{-25'd2305721}}, '{'{-25'd964211}}, '{'{25'd1551122}}, '{'{25'd628833}}, '{'{-25'd1634966}}, '{'{25'd964211}}, '{'{-25'd2054188}}, '{'{25'd2221877}}, '{'{25'd1718810}}, '{'{-25'd2557255}}, '{'{25'd2305721}}, '{'{-25'd1006133}}, '{'{25'd335378}}, '{'{-25'd964211}}, '{'{25'd1173822}}, '{'{25'd251533}}, '{'{-25'd377300}}, '{'{25'd2431488}}, '{'{-25'd1634966}}, '{'{25'd1593044}}, '{'{-25'd1173822}}, '{'{-25'd838444}}, '{'{25'd1718810}}, '{'{25'd880366}}, '{'{-25'd1089977}}, '{'{-25'd419222}}, '{'{-25'd1970344}}, '{'{25'd503066}}, '{'{25'd2347643}}, '{'{-25'd838444}}, '{'{-25'd2138032}}, '{'{-25'd2012266}}, '{'{25'd2389566}}, '{'{-25'd2976477}}, '{'{25'd1006133}}, '{'{25'd2557255}}, '{'{25'd1718810}}, '{'{25'd2389566}}, '{'{25'd377300}}, '{'{-25'd1425355}}, '{'{-25'd1593044}}, '{'{25'd1718810}}, '{'{-25'd544989}}, '{'{25'd586911}}, '{'{25'd670755}}, '{'{25'd1425355}}, '{'{25'd5324120}}, '{'{25'd419222}}, '{'{25'd2431488}}, '{'{-25'd1634966}}, '{'{25'd83844}}, '{'{-25'd1257666}}, '{'{-25'd754600}}, '{'{25'd586911}}, '{'{-25'd1593044}}, '{'{-25'd3102243}}, '{'{-25'd1341511}}}
};
