localparam bit signed [0:15][7:0] Output5 = '{-102, -30, -119, 33, -49, -93, -79, 37, 8, 89, 10, 124, -82, -73, 9, -58};
