localparam bit signed [0:46][15:0] Input4 = '{-16'd6983, 16'd13263, -16'd32393, -16'd16732, 16'd20329, -16'd21826, -16'd508, -16'd15887, 16'd24050, -16'd9011, -16'd23138, -16'd2707, -16'd2217, 16'd8930, -16'd28253, 16'd6729, -16'd29478, 16'd10167, 16'd1562, 16'd30070, -16'd3050, -16'd7732, -16'd1329, 16'd32098, -16'd4518, 16'd19507, -16'd1050, 16'd18222, -16'd16688, 16'd32317, 16'd26044, 16'd23343, 16'd30714, 16'd14440, -16'd28032, -16'd29302, -16'd12341, 16'd22413, 16'd28999, -16'd28066, 16'd5638, 16'd7853, 16'd15605, -16'd27234, 16'd13839, 16'd14505, 16'd6310};
