localparam bit signed [0:15][7:0] Output6 = '{-14, -14, -82, -38, 54, 109, -117, 40, 121, 69, -18, -108, -67, -87, -39, -20};
