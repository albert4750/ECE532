wire signed [7:0] convolve3_weight[4][8][3][3];
assign convolve3_weight = '{'{'{'{-24, 51, -90}, '{-39, -54, 115}, '{98, -5, -41}}, '{'{-32, -45, -102}, '{78, -96, -13}, '{70, -31, 44}}, '{'{-69, -71, 50}, '{45, 105, 4}, '{57, -35, -37}}, '{'{17, 35, 66}, '{20, 45, 57}, '{79, -9, 36}}, '{'{-23, 62, -124}, '{113, 114, 77}, '{30, -19, -41}}, '{'{98, 35, -55}, '{90, 55, -102}, '{-10, -106, 76}}, '{'{79, -30, -38}, '{-77, 102, -82}, '{80, -67, 60}}, '{'{-81, 122, -24}, '{0, 10, 75}, '{13, -57, -34}}}, '{'{'{-122, 45, 117}, '{30, -113, 41}, '{38, -75, 43}}, '{'{-46, 7, 92}, '{-63, 41, -62}, '{-14, -36, -50}}, '{'{101, 91, 118}, '{-28, 31, 93}, '{50, 124, 46}}, '{'{-35, -14, 33}, '{-116, 96, 105}, '{-48, -62, 72}}, '{'{115, -3, 10}, '{-16, 90, 27}, '{56, -8, -63}}, '{'{64, 69, -40}, '{-94, 79, -125}, '{60, 110, 37}}, '{'{43, 83, -40}, '{-58, 20, 6}, '{-100, -13, 6}}, '{'{-62, -36, 92}, '{-26, -27, -5}, '{69, -19, -55}}}, '{'{'{-28, 54, -51}, '{21, 123, 31}, '{-47, -93, 109}}, '{'{115, 122, 8}, '{126, -103, -107}, '{45, 101, 86}}, '{'{16, 25, 110}, '{-9, 37, -1}, '{1, 5, 70}}, '{'{12, -38, -54}, '{123, 54, -50}, '{-66, -56, 71}}, '{'{-83, 5, -81}, '{59, 42, 67}, '{10, 114, -71}}, '{'{91, -39, 3}, '{-3, 78, -46}, '{69, 58, 4}}, '{'{-111, 69, 63}, '{-34, 24, 3}, '{-59, 40, 36}}, '{'{-70, 49, 55}, '{24, 33, 18}, '{-31, 78, 113}}}, '{'{'{7, 53, 107}, '{-82, 112, 116}, '{-1, 33, -47}}, '{'{29, -116, -10}, '{-82, -10, -96}, '{-94, -13, -41}}, '{'{-4, 25, 46}, '{114, -21, -76}, '{105, -18, -64}}, '{'{-52, -10, -55}, '{18, -124, -121}, '{3, -80, -52}}, '{'{-91, -12, 109}, '{-80, -19, 82}, '{51, -79, -57}}, '{'{-38, 49, 110}, '{-99, -125, -54}, '{-44, 106, -63}}, '{'{-9, -108, 80}, '{-86, 114, -100}, '{26, -41, 52}}, '{'{-80, 66, -26}, '{-119, -126, -12}, '{-20, 105, -39}}}};
