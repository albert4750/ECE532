localparam bit signed [0:46][15:0] Input8 = '{16'd32240, -16'd1036, 16'd10879, -16'd1119, 16'd8529, 16'd21661, -16'd4596, 16'd28278, 16'd10030, 16'd27510, -16'd3808, 16'd7970, 16'd16499, -16'd27049, -16'd5508, -16'd3687, -16'd4946, -16'd22030, 16'd24427, -16'd460, 16'd24553, -16'd19858, 16'd5696, -16'd29364, 16'd28534, -16'd21943, 16'd4242, 16'd19204, 16'd18183, 16'd2691, 16'd9264, -16'd5044, -16'd26331, -16'd20364, 16'd9709, -16'd22992, 16'd6253, -16'd22574, -16'd22349, 16'd10801, 16'd11335, 16'd16218, 16'd11697, -16'd12306, 16'd5405, 16'd20995, -16'd24502};
