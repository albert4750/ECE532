logic signed [15:0] layer1_weight[20][3][9][9] = '{
    '{
        '{'{-30036, 10799, 9845, 19648, 13123, -11525, -2365, -665, 9225}, '{24275, -12011, 22258, 14116, -17833, -17338, 15832, 6744, 19852}, '{-18118, -15679, -538, -13785, 10327, 18606, -8616, 2897, 26277}, '{-15847, -5299, 6216, -25847, 6036, -30605, -27696, 4851, -24891}, '{-14338, -30897, -25169, -30272, 15186, -8093, 10200, -847, 755}, '{-31971, 17043, -29549, -17522, -7769, 23840, -16447, 19721, -13639}, '{21119, 8736, 23071, 17098, -14092, 24727, 27299, -1538, -21045}, '{11122, -15177, 22556, 25378, 10368, -6016, 26532, -9163, -26747}, '{-12762, -29208, -7436, 28945, -1713, 12676, 18025, 27690, 13754}},
        '{'{14879, -11400, -12031, 30017, -4121, 28585, -6087, -18141, -20634}, '{27767, 15115, 8622, 23634, -12197, 30592, 27022, 19043, -22987}, '{-13428, -5511, -16470, -20396, 18635, -28348, 13062, 7108, -15313}, '{29311, -18444, 5251, 29644, -25756, -23372, 14312, -28850, -23409}, '{18068, 11491, -9286, -17641, 10959, 2957, 4469, -18603, -24016}, '{30001, 9797, -18263, -26973, 17856, -9121, 7365, -4514, 8448}, '{22385, 3762, 29988, 26530, -7376, -16547, -13949, 1634, 15914}, '{-31795, -11920, -22553, -21611, -7991, 27007, -18944, 30602, -30350}, '{-19925, -19526, 3455, 22551, 22203, 28802, -26247, -10142, 24126}},
        '{'{-23645, -1314, 30843, 10179, 23122, -18514, 19171, -9068, 4305}, '{18994, 5531, -9458, -983, 31802, -17727, 23588, -9462, 4182}, '{15403, -19608, -6133, 15106, 307, -19376, -18400, -27466, 1152}, '{-9434, 8467, 5294, 13866, 13683, 17592, 2492, -5656, 15949}, '{14622, -19176, -7555, 770, -16893, -24482, 11490, 5995, 32013}, '{30576, -14040, -19128, -29677, 12895, -28856, 17818, -26174, -11016}, '{24756, 26947, -9236, -24771, 20238, 8032, -17148, 8131, -27923}, '{-6005, 21500, 10838, -29235, -29831, -6547, 4939, 31416, 9744}, '{-13160, -27747, -5995, 1134, 16409, 9680, -15428, -30855, 19318}}
    },
    '{
        '{'{-19339, 26045, -18861, 2721, -22680, 17312, -17180, 5627, 27387}, '{22649, 5446, -32299, 10527, -24051, 18247, 1720, 5272, -15793}, '{6185, 18706, -16856, -4682, -16177, -17653, 20646, -18321, 19805}, '{-4103, 21633, 31455, 10102, -21716, 24792, -17027, 24600, -4029}, '{11218, -27665, 24323, 2282, -31028, 22502, -20189, -26922, 13310}, '{15037, -12603, -29993, -13781, -2016, -9205, -18840, -26412, 1162}, '{14006, -4117, 30117, -16771, 32412, 623, -536, -23806, 30235}, '{-12333, 1241, 10903, 25397, -28365, -15186, -2924, -13387, 5661}, '{-16829, -21981, -15577, 28041, -30647, 12585, 31639, -8317, -28882}},
        '{'{8922, -10318, -17556, -22781, 18207, 15113, 28042, 28187, 12717}, '{-16185, 1447, -27587, 10581, 29537, 27692, -21726, 10146, -27560}, '{-26591, 14981, 30952, -27905, 22564, 18176, 17867, 14626, -24379}, '{-31874, 30645, 21758, 15440, -2626, 136, -5955, 6273, 26833}, '{-6800, 14627, -19080, -29349, -16216, -26764, 2852, 12464, 9753}, '{-11965, 24423, 25084, -17629, 3186, -10466, -11235, -14607, 19745}, '{8338, 21777, 20701, -18092, -11779, -30206, -10171, 30053, -7284}, '{4652, -19595, -5379, 13634, -4497, 22619, -21163, 423, 28199}, '{32715, -4458, 28062, 28305, 23238, 967, 4370, 9052, -10197}},
        '{'{21587, 433, -19671, -10147, 29870, -14955, 28873, 12121, -13838}, '{-1568, -18469, -16055, -12772, -16405, -7983, 23145, 30650, 3968}, '{-8234, -449, -31728, -26518, 24740, -7586, -25064, -25996, 5311}, '{9411, -6861, 12424, -23624, 29531, -5027, 6011, 19182, 29783}, '{8352, -30573, -28088, 22983, -7081, 19469, -710, 22097, 5240}, '{-22668, 27575, -17600, 10955, 732, 21412, 24857, 13088, -8790}, '{-20722, -11818, -23268, 7444, -46, 19780, 13846, 21731, -9350}, '{16979, 647, -20536, -15811, 6797, 5637, 24832, -4984, 11471}, '{14799, -75, 5259, 9220, 6567, 4444, 19373, 29978, 586}}
    },
    '{
        '{'{-18636, 21486, -25167, -4901, -21709, -32029, -3223, -11502, -4747}, '{-27358, 15923, 16030, -15947, -28870, -4181, -14537, -23044, 17404}, '{-9454, -31827, -5289, -7743, -21178, 21994, -21451, -23760, -930}, '{-14277, -18096, -6502, -2436, -12125, -20934, -15439, 29802, -24375}, '{23852, -14579, 15225, -30906, 8742, 3751, 9864, 31757, 18424}, '{-31865, -2352, -17416, 31254, -7688, -8369, -18471, -26872, -20765}, '{-24826, -9007, 9671, 31188, 5593, -16446, -2500, 29072, 19512}, '{7026, 3821, -13673, -24296, -31740, 2660, 29676, -30415, -5801}, '{-10722, -25034, -8039, -4332, -8863, -5787, -21831, 12695, -613}},
        '{'{-31715, -13407, -10893, 3893, -30089, -21581, -27818, -1546, 28679}, '{-30103, -13327, -1911, 6838, 3968, -31917, 25976, -27740, -12591}, '{-9068, 24437, 7152, 19715, -8066, 22314, -23999, -10732, 804}, '{5444, 19408, -16272, 1967, -15734, 4333, -31384, 13278, 30555}, '{-18901, -32705, 3999, -28780, 18886, 29961, 19900, 12891, -13713}, '{13731, 2387, -6324, -10990, 3441, -24758, 26850, -19231, 18347}, '{-27005, -13428, -25372, 3898, 20353, -18063, 23680, -11481, 29720}, '{-7494, -16092, -1693, 25413, 14470, 20483, -27422, -9351, 4776}, '{-1604, -19039, -8932, 23364, -28646, -32032, -5896, 4461, -14413}},
        '{'{-21303, -19019, 8389, 13217, 1671, 27261, 606, -14264, 12534}, '{23380, 25735, 18115, 26837, -16933, -24980, 19779, 6246, -8364}, '{-5817, -7597, 5343, -30464, -20859, 3419, 1131, -1122, -18487}, '{-14381, 28167, 27797, 10213, -8740, -19064, 18091, -22994, -24576}, '{-25240, 691, 13862, 29785, -5046, -13837, -5406, -30085, -7849}, '{-17312, -25773, -3814, 23246, -26592, -5005, 6598, -26783, 4524}, '{827, -22727, 23218, -22355, -2327, -29564, 28089, -32675, 15707}, '{-19055, 2467, 3778, -32364, -27731, -6983, 13263, -32393, -16732}, '{20329, -21826, -508, -15887, 24050, -9011, -23138, -2707, -2217}}
    },
    '{
        '{'{8930, -28253, 6729, -29478, 10167, 1562, 30070, -3050, -7732}, '{-1329, 32098, -4518, 19507, -1050, 18222, -16688, 32317, 26044}, '{23343, 30714, 14440, -28032, -29302, -12341, 22413, 28999, -28066}, '{5638, 7853, 15605, -27234, 13839, 14505, 6310, 13621, -29781}, '{-11694, -4729, -29476, 19265, 5801, 31554, 23666, -21668, 8526}, '{-7451, -6949, -778, -24476, 18847, -22307, 29874, 7676, -8018}, '{-7587, -24974, -12639, 4876, -12576, 9961, 9040, 25666, -10808}, '{-3085, -30595, -23414, -11664, -25894, -15205, -7496, -9096, 28993}, '{-13888, -30011, -20648, -8926, -28721, -14333, 23228, 19694, -24923}},
        '{'{31915, 18131, 11096, 32326, -24940, -7290, 3868, -11661, 4998}, '{-27838, 16988, 24540, 3686, -7323, -12933, -12603, -19347, 9545}, '{-32668, 21174, -23731, -26731, 22011, -7521, 20049, 19491, -7955}, '{15603, 14586, -1656, 23294, 9497, -16363, -9811, 17637, 6102}, '{-7792, -2919, 25582, -29577, 9893, 8063, 30081, 30085, 18118}, '{6540, -29350, -23990, -1029, 21430, 7246, 9022, 26184, -1849}, '{32557, -13179, 15919, 29371, -11094, 20931, -26486, 21234, -31431}, '{3547, -19111, -15997, -27523, -5426, -28846, -31547, 14010, -30844}, '{23569, -23867, 8639, 16734, -23912, -12669, -3771, -24152, 4260}},
        '{'{24122, 9393, -29257, -21864, -32095, 1938, 24417, 12750, -7439}, '{-25465, 18357, -3349, 28718, 32240, -1036, 10879, -1119, 8529}, '{21661, -4596, 28278, 10030, 27510, -3808, 7970, 16499, -27049}, '{-5508, -3687, -4946, -22030, 24427, -460, 24553, -19858, 5696}, '{-29364, 28534, -21943, 4242, 19204, 18183, 2691, 9264, -5044}, '{-26331, -20364, 9709, -22992, 6253, -22574, -22349, 10801, 11335}, '{16218, 11697, -12306, 5405, 20995, -24502, -428, -9750, 11585}, '{6007, -29164, -29488, -27606, 5618, 16412, 1434, 2903, 3252}, '{-26320, 14274, -6554, -7415, -25342, -21132, 31596, -2327, 13145}}
    },
    '{
        '{'{13692, -7307, -32156, -28582, -7100, 25193, 9738, -12276, 22120}, '{10465, -5723, -12121, -23648, 25978, 11553, -23654, -32669, 23769}, '{-30414, 26968, 31954, 22292, 13022, 32412, -31160, 21778, -2663}, '{-7272, -25049, -21270, -18821, 16668, -2408, -20846, 32451, 14508}, '{16083, 26925, 11062, -16384, 26762, 21187, 30598, 5851, 14179}, '{10681, 28614, 19347, 25762, -30670, 14578, 4966, -30700, -25941}, '{-19850, 26752, 5604, -9875, -20375, 7874, 24801, -8564, 1807}, '{-13194, -17887, -5993, 1932, 3973, -986, 28417, -32502, 11270}, '{-131, -27386, 8806, -4186, 12619, 30066, 25941, -4738, -13966}},
        '{'{-9550, -205, -4862, -25268, 4765, 22025, -23949, -7224, -28283}, '{-9612, 24757, 2283, 20673, 32555, -1457, -21442, -5812, 14895}, '{-9652, -2411, 16504, -18670, 14681, -7667, 16606, 3676, 20716}, '{-22423, -21291, 11782, 12900, -12752, -6616, 9114, -25442, -25211}, '{14479, 13247, -21019, 11301, -453, -16783, -20385, 14688, 2544}, '{14544, -26336, 62, -5750, 27020, -2467, -16576, -2659, 6490}, '{-30745, -24426, 24979, -13947, 2852, -3501, 16511, 1508, 9989}, '{-17060, 18892, 23706, 12017, -7085, 12172, 2022, -7033, -13132}, '{-32176, -9827, -15360, -12585, -1329, 32586, 32508, 28291, 4669}},
        '{'{18755, -21360, -22672, 9673, 7764, 116, 25317, 7935, 824}, '{30014, 23480, -9680, -11119, 26485, 8121, 3593, 12780, 21694}, '{-6065, 25318, 23758, -7775, 26500, -5232, 2276, -30905, 23870}, '{16151, 32603, 26990, -24569, 6653, 8982, 1890, -5986, 26358}, '{1616, 25755, -16849, 20975, 626, -17909, 22487, 22350, -20505}, '{-7394, -30630, -1758, -5578, -6319, -9565, 23623, 7021, 16187}, '{-19856, 4517, -3004, -24139, -5107, 22629, -3309, 32619, 11528}, '{-25760, -14639, -2875, -5764, -24476, -31359, 765, -11107, -27771}, '{-8240, 20710, 12792, -26712, -30058, -13282, -18177, -9709, 9988}}
    },
    '{
        '{'{21140, -25750, -13750, 123, 15811, -810, 6460, 27365, -2822}, '{-14755, -3415, -27096, 26812, -23343, -3405, 1320, 14395, 2538}, '{-23074, 18973, 14561, 7774, 23790, 11941, 20862, 10456, -752}, '{-25757, 23719, 7837, 25084, -13247, -16617, 27848, 1408, 1111}, '{3877, -10897, -5697, -5734, 21209, -19111, 15494, 14552, 17911}, '{27087, -7067, -15063, 26513, 32720, 3952, 3115, -15250, 19909}, '{20854, -29805, -9489, 14102, 28013, 8075, 31243, -17503, -8313}, '{-6025, -28390, -7632, -21305, 12527, -13642, 21088, -28316, -6318}, '{-26025, 9621, -27138, 18946, 11528, 23818, -5883, 3366, -25690}},
        '{'{-23964, -11839, 26229, 571, -12636, 17285, 18693, 6182, 11939}, '{-10152, -16463, 5839, -684, -9870, -23287, 12279, 7300, 31665}, '{-13288, -22946, 19842, 24403, 20355, -12723, -31477, 24973, 2532}, '{2129, -7014, -20538, 18095, -2462, 30229, -20588, -26966, -24710}, '{18873, -15215, -3483, -12327, -4876, 6613, 16567, -16796, -4924}, '{-28561, 21730, 19211, 12258, -26527, -14098, -1645, -16528, -11253}, '{7137, 13849, 5217, -27297, 18733, 19206, -17831, -20648, -5651}, '{-30170, 4147, 9232, 24471, 28378, 21251, 1882, 12718, -24966}, '{21917, -3326, -32123, 21881, -28729, 23311, -9394, -23133, -10060}},
        '{'{-10905, 16246, -9977, 10931, -21146, -32007, -23629, -12387, 4791}, '{625, 8587, 27075, 5837, -20614, 3383, 32344, -30213, -17156}, '{20984, -2236, 27765, -18061, -554, -27463, -1699, 6758, -19573}, '{16078, -25006, 28633, 3308, -4093, 165, 1415, 18205, 9294}, '{28427, -21559, 16907, -1264, -25540, 27259, 24679, 14015, 699}, '{-10111, -18542, -20811, -19172, -15936, 29525, -20776, -2487, 15240}, '{-8238, -29301, -22052, -9867, 14259, 27473, -3657, -29681, -32637}, '{29802, 27096, 16597, 3356, -4294, -20779, -31154, 2927, -7359}, '{4940, -31477, -6887, -15001, 30475, 25434, -27923, -10846, 30593}}
    },
    '{
        '{'{19454, 17040, 11521, -22000, -30175, 19489, 23724, 1510, 9000}, '{-5816, 26829, -31638, 595, -27918, 17824, -11369, 16708, -27233}, '{8854, -9152, 7909, 32031, 79, 24659, 23311, 11059, 32249}, '{11660, -5459, -27638, 22004, 9833, 9040, -5050, 30741, 11998}, '{-31037, 17744, -10944, 9345, -6350, -17568, -16021, 29691, -28206}, '{18770, -23879, -12906, 7951, -23665, 11804, -29369, -19173, -18216}, '{-28359, 19258, 10456, -2100, -14067, -26734, 16462, -24626, 22292}, '{-27065, -2377, -4820, -1813, -8971, 19547, -10196, -24817, 10237}, '{-14761, -26677, 1613, 8702, -25187, -10657, -3986, -16686, 7812}},
        '{'{-3556, 30401, -6095, -27727, -13993, 15929, 7888, -25559, -23078}, '{18160, 9410, 7087, 18705, 31764, -1370, -31424, 32390, -16148}, '{-3434, 18511, 6218, -15198, 28328, 6822, 19446, -10603, -8414}, '{8565, 11424, 18858, -6785, 15660, -32157, 30505, -9479, 15207}, '{-28773, 14075, -30416, 21887, -14710, 13636, -23279, -9469, 24165}, '{22110, 29143, -22243, -19866, 1659, 7326, -11061, -3646, 19933}, '{-25284, -5497, 6835, -26380, 10825, 11735, -18496, 30704, -3695}, '{13992, -16141, 2581, -2466, 14234, 3215, 2800, 14097, -9974}, '{-14703, -18301, 19431, -439, -15587, -9021, 27079, 4560, 2274}},
        '{'{-20860, -7747, -2214, -7068, 14470, 28704, 11345, -14729, -30346}, '{18165, -26331, 14967, -15077, 29747, 13902, 16315, 5718, -31137}, '{-6136, -13000, -9443, -1380, 18399, 21922, -24390, 22399, -28802}, '{-12335, -27172, 26735, -8560, -4152, -10693, 12535, -31764, -11257}, '{-5236, 13600, 20180, -11541, 28747, -29475, -31704, -19456, 24788}, '{25709, 14940, -819, -19291, 31151, 29245, 4199, -2126, 25156}, '{-24082, -25652, 16057, 9079, 12261, -28688, -19324, -1431, 2596}, '{29008, -22062, 16549, -23842, -16011, 26094, -8925, -10320, 13952}, '{22065, -13127, 20745, -10190, -5407, 9392, 24561, 29196, -4410}}
    },
    '{
        '{'{15996, -13837, -18524, 13411, -3738, -11228, 23838, 22130, 23699}, '{-4698, 29100, -16349, -11506, 22557, 16307, 16444, -19464, -25263}, '{23363, 26397, -20325, 15491, 17441, 32501, -11853, -28810, 1435}, '{3300, -24520, -26347, -3417, -12566, 7498, -13795, -5903, -5219}, '{957, 9786, -26856, -12174, 11536, -26176, -12444, 30690, -17797}, '{-6131, 769, 28411, -28414, 1858, 10387, -22028, -12550, -27188}, '{-29026, 1575, -555, 5709, 2993, 1306, 12659, 17548, -29455}, '{17344, -22271, -12892, -16630, 20330, 22816, -23042, -25316, 27322}, '{15042, 2780, 29761, 17613, 31059, 6703, -17839, -3676, -825}},
        '{'{-6859, 9926, -11639, 19983, -9454, -31587, 29365, 3004, 12842}, '{-30254, 23170, -21731, -18031, 18467, 31608, 3347, -12400, -12777}, '{-24948, 4451, -25747, 14008, 26306, -25836, 15491, -20399, -13396}, '{-30682, 23594, -9270, -19931, 362, -28120, 18287, -20709, -18812}, '{1459, 27030, 10917, 6947, 542, 18183, -25640, 13912, -32529}, '{-18545, -5750, -25453, 2893, 6119, 22328, -26651, 16359, 10130}, '{7623, 16444, 24600, -20320, -29332, -8921, -1164, 31848, 13694}, '{367, 4212, 26596, -18454, 20496, -19532, -10022, -20504, 26832}, '{25390, -25376, 2654, 18260, 20247, -12657, 20652, 14931, -27529}},
        '{'{-14793, -19102, -21093, -26323, 23522, -19119, -28969, 32155, 28237}, '{-32336, 26583, 11102, -10875, -7815, 20711, -3359, 17265, -19486}, '{18204, -4876, 15425, -14268, -1323, -5688, -26884, -32398, 7073}, '{-19082, 7651, 26160, -11165, 8153, 13893, -18495, 18019, 26695}, '{-5631, 16513, 4295, -20839, 9316, -13747, 7788, 3250, -31333}, '{-28576, 17963, -28909, -9886, -15059, -24476, -11952, 28784, 27882}, '{21369, 23467, 15811, 14856, 30931, 31662, -26048, -32396, 28564}, '{-29600, -14878, -3221, -1659, -20139, -26344, 9218, -9731, 31741}, '{3527, 29804, 2251, 243, -228, 16758, -19617, -28607, -30256}}
    },
    '{
        '{'{22898, 28882, 11662, 15893, -2961, -10385, 6341, -23775, 15978}, '{-11134, 12827, 27368, -11913, 15507, -28785, 4935, 18412, 6941}, '{17827, -13599, -18128, -31823, -31920, -3912, 16703, -25128, -6726}, '{-19579, -2253, 21754, 21053, 19562, 27091, 23825, -30675, 5088}, '{9790, 19478, 29921, -8602, 28297, 31493, 17740, 30269, -5974}, '{-15625, -11888, 3387, 28945, 31940, 17724, -26983, 5262, -31891}, '{-24771, -3915, -32687, 28189, 2246, -20452, 16074, -379, 31204}, '{-19996, 31060, 12215, -11790, -28494, -29098, -26443, -6390, -4565}, '{-21573, -6754, -26821, 9358, 26611, -19024, -11656, 30077, 1080}},
        '{'{-11839, 1896, -121, 31685, 10383, 8823, 3049, -22220, 6432}, '{11351, 14286, -29790, 22045, -10189, 24025, 8629, -5372, -27456}, '{3963, -14182, -6700, 2437, -1670, -25768, -30447, -22588, -30408}, '{-22368, -19215, -32431, -2488, 16457, -15644, -2657, 26974, -4791}, '{29036, 3248, -32029, -19040, 5390, -11715, -4777, 24992, 26936}, '{-24164, -28501, -19359, -16206, 27438, 26732, -10424, -13915, -5512}, '{10242, -23791, -12145, -15677, -23211, 22000, -3342, -13219, -18587}, '{15480, -17770, -27438, -8697, 9015, -22351, -11238, 29432, 25220}, '{-17299, 24665, 29722, -324, 10483, -12689, -10669, -17842, -28014}},
        '{'{11385, 19040, -22181, -5340, 32102, 32148, -6785, -27156, 24963}, '{18066, 8397, -6093, -3535, -481, -1567, 22162, 18700, -9617}, '{32731, 30951, -21662, -8377, -4514, 6957, 3792, -22463, -14248}, '{14608, -26323, 22911, 6363, 165, -15950, 14744, 1968, 1228}, '{-23548, 21488, -11341, 1198, 31784, -4210, 11505, -18038, -25189}, '{3406, -27802, 5517, 19972, -11562, 21775, 7197, -23602, -9046}, '{32409, -15157, 12767, -8997, 18966, -25490, -3285, 1492, 3767}, '{-17667, 17538, -8551, 26237, -1928, -14720, -12961, -32584, 7278}, '{11974, -27694, -1450, 10430, -257, 7726, -19717, 5209, 19149}}
    },
    '{
        '{'{18060, -26306, 16677, 20435, 14495, -27785, -24676, 26939, 30200}, '{-3757, -4312, 9576, -2695, -8615, -20497, -28899, 31516, -7116}, '{32042, -5494, 3796, -27375, 25216, 11943, 28710, 1506, -7999}, '{-16848, -18218, -25555, 1146, 2737, 30230, -3865, -10754, -17060}, '{-15039, -31403, 30530, -18912, -13902, 25926, 27238, 23459, -6155}, '{25060, -14185, -16397, -30598, 18514, 5222, -16295, 25326, 30799}, '{-29583, -24421, 24405, 1537, 2313, -20365, -30895, -20085, -11200}, '{2295, 5955, -12807, -835, -8138, -15068, 31188, -4994, -24557}, '{1007, -12603, 4820, 23165, -16706, -828, 21673, 16592, -13680}},
        '{'{2233, -16763, -6048, 2326, -2941, -14968, 21310, -6308, -31575}, '{10058, 24678, -22948, 15455, 18540, -31861, 21410, 16475, 18225}, '{12871, 26023, 27494, -17545, -966, 29701, 1097, 18264, 12428}, '{2792, 25825, 28475, -11570, 14317, 11791, -23548, 30614, -31052}, '{14402, -12473, -25235, -5816, 3333, 25127, -24241, 12111, -4311}, '{15321, 662, -17959, -23335, -11373, 7998, -23779, 9993, 28043}, '{-21635, -10141, -486, -21657, -2817, 3794, -25016, -16129, 30337}, '{-8349, 6770, 6385, 32430, 9527, 26122, -16694, 5400, -1537}, '{-10913, 29739, -3109, -31091, -11314, 20535, -26619, -7785, 22570}},
        '{'{-27033, -17359, 17765, -3226, 26187, -14475, 23480, 32171, -28520}, '{-12975, 30229, -10274, 19602, 12351, 21849, 1565, -8923, -13391}, '{-11096, -28175, -22166, 23775, 20583, 3339, 24888, 24565, 7615}, '{22670, -23264, 6337, -27527, -16011, -31935, 22564, -18694, -30695}, '{-20532, -26552, 30770, 14860, 2968, 12435, -2365, -9846, -9721}, '{-15436, -17316, -498, -13880, -4050, 5347, 12323, 2257, -31593}, '{10301, -10635, 17589, -11764, 5549, 32263, 29178, -10833, -22418}, '{-7513, 32606, 5779, 1258, 1901, -27726, -16831, 19371, 16978}, '{-14898, 30715, -2983, 101, -5768, 20664, -17848, 6834, 10274}}
    },
    '{
        '{'{17370, 8715, -13716, 3211, -22168, 6564, -12418, 19633, -12340}, '{22481, 21727, 20426, 5936, -11702, -4981, -17827, 5666, 13002}, '{3532, 2801, -25305, 26992, -6646, 25346, -6791, -27665, 75}, '{-30802, 19507, 23028, 12201, -28678, 31835, 3715, 18704, -17089}, '{-17600, 7949, -28890, -28412, -17917, 25491, 21073, -29552, -30338}, '{31559, 8856, 9483, -8042, -12740, 9435, 21122, -27768, 21576}, '{-2343, 6438, -31180, -287, 18776, 15679, -21611, 31236, 18847}, '{-23821, 14539, -1371, -2297, -12650, 28284, -6870, 22715, -21793}, '{16694, -10295, -16525, -19021, -5550, -4329, -17325, -10471, -10439}},
        '{'{23749, 22873, 16685, 15727, -2472, -6221, -31429, -14420, -15206}, '{3704, 19061, 31659, 21113, -7776, -6370, -26994, -12985, 28768}, '{-14659, 513, 3574, -18001, -25220, 18797, 11382, -9045, -13862}, '{25615, 8004, -15158, -10155, -4441, 106, -25109, 13918, 32214}, '{-28416, 9809, 19642, -5108, 21723, -17621, -27722, -1667, -7761}, '{-23786, 15135, -20108, 15394, 26594, 28458, -29372, 3962, 17214}, '{3876, -4269, -5972, -23855, -22288, -17041, 8390, -7930, -29264}, '{30089, 24092, 20557, 30392, -30327, 469, 26434, 14857, 29806}, '{7160, -31580, 8476, 22004, -17344, -15414, 13180, -2931, -789}},
        '{'{26114, -30299, -9273, 7255, 1758, 4049, 26115, -16273, -18462}, '{-25776, -30989, -28078, -11470, 18365, -30230, 29650, -20452, 1827}, '{24885, 12058, -29327, -27289, -27094, 28462, -3899, 23068, -8065}, '{24747, -23469, 20542, -1206, 11466, 23177, -15141, -27933, 15179}, '{-13472, 28838, 22559, -20749, -8298, -29314, -2213, 5945, 23573}, '{28385, -28867, -532, 3881, -1677, -11413, 26979, 31913, -5894}, '{-24937, -8963, -29976, 5940, -32489, -23430, 20296, -20951, 19693}, '{-19652, -31953, 9871, 29732, -26687, 2654, -22555, -15574, -8450}, '{512, -45, 19334, -27939, 3139, -28385, -29923, -26608, -6205}}
    },
    '{
        '{'{-1766, -12291, 25862, -12055, 11749, -12021, -29359, -21705, 4989}, '{-23253, 6467, -19948, 12763, -32257, 19063, 13788, -28402, -16114}, '{-6064, 15843, -32321, 4469, 16102, 43, 31899, 7526, 11991}, '{5012, 29691, 2583, 5410, 3360, -29887, 29974, -29931, 29113}, '{19012, -8403, 1000, 28583, -11496, 10582, -18159, -12364, 28122}, '{3720, -5371, -11039, 12630, 24826, -20910, 22282, 2622, 1565}, '{139, -22370, 8519, 3642, -19490, -2006, -8235, -9913, -7527}, '{492, 17206, 21622, -16045, -2023, 26797, 1401, 16874, -25469}, '{-31884, 7124, -28687, -31917, -14087, -30171, 30881, -9796, 17260}},
        '{'{11993, 26119, 19388, -1883, -16812, 23546, 20834, -1776, 13997}, '{-31256, 23719, 7713, -8351, -6335, 22729, -10153, 5444, 14616}, '{-7162, 24417, 1394, 21247, -20932, -808, -14275, -9228, -9029}, '{19959, 15993, 10698, -11491, -31505, 25592, 4124, -9064, -4733}, '{4562, 26261, -13050, 14420, 17685, -29065, 32027, 2970, 8153}, '{29120, -1682, 27011, 30517, -25819, -18425, 1400, 15696, 7627}, '{19083, -6164, 14722, 7478, -23035, 27409, 24314, 8061, -25010}, '{-18555, 31566, -19375, 9449, -32658, 2668, -31714, 20322, -22781}, '{-32640, -14499, -22228, 31404, -15124, -12417, -5517, -5187, 18686}},
        '{'{3072, 28433, 18845, 18011, -19550, -31758, 23539, -23324, 1211}, '{-19435, 12351, 22238, 15864, 26213, -17775, 23590, 9935, -21631}, '{-18289, -5143, 6870, 18157, -8687, -15124, 10165, -17002, -18995}, '{2674, -4945, -6462, 24843, -30839, 31218, 27432, 12214, -31821}, '{-4049, -7420, 30602, 11761, -18178, 29318, 11638, 19884, 15688}, '{32136, -10040, -15892, 12005, 12306, 29698, 10437, -17187, -15879}, '{17637, 30308, 362, -30563, 9371, -9583, -3654, 16779, -29391}, '{-19128, -28328, 26115, 18032, 30731, 20281, 3506, -16753, -4167}, '{16515, -8330, 23524, -26692, 10151, -18946, 26581, 20637, -13387}}
    },
    '{
        '{'{12355, 9784, 22731, 23927, -11185, -5843, -28070, 2127, 23777}, '{-11253, 7671, 26757, -15458, -4934, 1604, -7877, 8736, 20261}, '{7339, -23939, -17092, 12845, -26339, -16134, -23397, -4377, 17179}, '{29725, -24450, 6216, -27573, 26721, -29490, -4570, -21237, -29238}, '{18166, -24743, 22560, -22862, -25560, 9414, -26338, -14698, -23429}, '{-12725, -2781, -28204, -13372, 9791, -27900, -3407, 4980, 9373}, '{22207, -17603, -32165, -401, -9005, 24936, 6234, 11802, 25161}, '{6066, -22305, -12450, 10001, 26311, -24776, -17421, -1245, -24375}, '{26332, -20689, -30672, 29047, -13369, -9611, -5565, 20091, -8505}},
        '{'{2366, -17464, 18725, -29691, 7777, -32713, -25124, -2642, -30682}, '{-19919, -30456, -390, -6975, 5442, 21566, 26640, -11075, 28866}, '{-17141, 22943, -29302, 4116, 9316, 5902, -29064, -32716, 8647}, '{-16739, 18309, -13042, -22926, -15634, 27599, -31949, -25568, -7785}, '{-10503, 25435, -27898, 30409, 26744, -3007, -31669, 25431, -30212}, '{-26938, 11048, 28348, 21540, 13196, -11357, -8130, 1477, 30526}, '{-32326, -11700, 28178, 10624, 1025, -18732, -15667, -22950, 13424}, '{-917, 13461, 30286, 29965, 5096, 19523, -14487, 22929, 30981}, '{-16358, 31423, -2661, -21, -22803, 32681, 21005, 31533, 28080}},
        '{'{-24008, -24518, -5103, -2858, -17569, 31705, 6364, -819, -7801}, '{10522, 6417, -25916, 22059, -5713, 11998, 22653, -15012, -12807}, '{-24760, -12614, -24805, 10246, 903, 2741, -20617, -18952, -22502}, '{3707, 21195, 16165, 17501, -11855, -16876, 20957, -13449, -26184}, '{-8259, -3657, 29404, 24727, 19129, 22153, -30080, -410, -15981}, '{14791, -13262, 31270, 31683, 30460, 3486, -29147, 22456, -30850}, '{4073, -19835, 12347, -24624, 21978, -11843, -2273, -31802, 31065}, '{-29493, 9873, 19487, -11617, 20564, -12198, -3033, 757, 18610}, '{17994, 14630, 6724, -22149, 12839, -28545, -21297, 16397, 25763}}
    },
    '{
        '{'{8678, 26491, -12917, -32409, -11957, 22512, -18634, -2652, 5202}, '{-5941, -13645, -26462, 22458, 80, 540, 14729, 30565, -4088}, '{12433, 30448, -7956, -6948, -6503, -29346, 11387, 101, 5819}, '{25979, 24542, -11271, -3013, 9402, 3346, -26100, -29823, -19173}, '{21002, -22589, -22595, 784, -741, 19068, 3846, -9728, -10233}, '{31385, 22595, 1851, 20216, -9868, 12799, 6564, 14764, 3797}, '{31345, -14602, -1537, -13112, -1425, 19622, 1962, -13343, 24228}, '{-10172, 28763, 8973, -371, 11177, -16056, -9594, -23202, -7028}, '{8802, -14461, -5912, -25072, -30459, 20008, 9655, 15261, -14667}},
        '{'{-7914, 29029, -13801, -24325, -28806, -23644, -8469, 12475, 11298}, '{7110, -9850, 344, 26188, 5137, 30303, 9776, 20261, 15360}, '{3530, -25999, -5268, -25596, -8609, 25532, 1663, -9718, -27875}, '{29537, -10391, 1264, -31219, 4371, 16425, 29900, 7596, 14387}, '{-7061, 26768, 19960, -4098, 10994, -28763, 9742, -15708, 15474}, '{-19324, 8178, 303, 10112, -20687, 19365, 28926, -20021, -9428}, '{-10683, 24936, -15890, 26384, -2800, 18186, 3589, -25705, -9297}, '{-6589, 7334, 7152, 10514, -26530, 24016, 14111, 31146, 30767}, '{7445, 5089, 19511, 1354, -22420, -7137, -15789, -958, 4243}},
        '{'{-21345, 32626, -13549, 2855, 22439, -1475, -32159, -20564, -22284}, '{-20756, 16822, -20770, 25722, -17945, -26434, -26420, 13200, 80}, '{-30210, -23418, -2620, -11475, 15316, -9734, 9886, 12876, -22661}, '{-27979, -4703, 602, -27246, 19590, -23944, 5250, -13158, -26386}, '{-20199, 27149, -2113, -13605, -13762, -13255, 2341, 21421, -29291}, '{-32661, -24072, -27835, 5113, 26417, 5145, 16652, 15924, 19270}, '{31663, 8957, -32695, -21622, 6728, -28198, 21648, -31393, 8030}, '{4862, -29467, 2342, -15184, -14660, 16902, -5136, 13254, 17015}, '{-7679, -18065, -23361, -4927, 26237, -15083, 814, 9984, -20778}}
    },
    '{
        '{'{-13148, -20838, -14700, -20140, -25369, -27102, 30961, -21650, -5059}, '{18334, 27291, -13596, 1609, 11592, 22068, 15956, 17303, 28990}, '{-4048, -6169, -2629, -23253, -24662, 653, -32264, -32401, 9209}, '{-7415, 19611, 32346, -31771, -2526, 5958, -19031, 32749, 13349}, '{12294, -4806, -11691, -27645, -18357, -12566, -4853, 27037, 6222}, '{-11565, 5402, -1685, -25857, -12208, 25763, 1588, 5009, -432}, '{22922, 24569, -27460, -31799, -20381, -19559, 18047, 19610, -15821}, '{-24241, 18715, 26756, 19814, 24277, -6041, -30479, -22091, 3863}, '{5100, 16358, -25237, 6763, -14826, 1372, -28690, 7211, -3066}},
        '{'{-31859, 17613, -3951, 7592, -25987, -24098, -10812, -22766, 8944}, '{-27518, -16357, 16776, -28949, 21711, 5683, -32553, 30639, -21697}, '{-13154, 14861, 11100, -1106, -4210, -24846, -850, -4947, 22113}, '{-3836, 21364, -28022, 30068, -8129, 12562, 3556, -14136, -28553}, '{-14022, -20791, 15086, -29299, 7692, -19811, -13746, -9880, -32691}, '{24201, 28590, -27972, 588, 13541, 28317, -17299, 28747, -16916}, '{-6167, 10097, 26520, 12091, 32712, 6799, -17994, 4768, 25068}, '{-11010, 11984, 5106, -26253, 28268, 9330, -17039, 12299, 2319}, '{13593, 21269, -14186, -18479, 31708, 17146, -14501, -3988, 29128}},
        '{'{-31909, -20004, 27367, -17813, -3993, -8093, 22942, 5876, -87}, '{-26890, 12681, 17270, -7372, -4821, 27473, -2126, -10864, -960}, '{-22758, -18297, -23114, 15186, -70, -15029, 6457, -8518, 27596}, '{10509, -15416, 232, 7954, 27793, 29866, -13012, -13086, 9931}, '{27479, -19642, -1842, 11822, -16842, -8526, -32725, 8769, -5170}, '{-20123, -18170, -14215, -2897, -29524, 19209, 515, 25993, 28795}, '{32500, -22021, -11230, 19934, 23041, -27354, 26830, 6096, 19294}, '{11698, -24435, 5974, 30766, -1053, -23721, -23771, 12125, -20755}, '{31466, 19802, 24658, 4054, -28154, -6582, 23979, 18945, 3529}}
    },
    '{
        '{'{14810, -28496, 6991, 13713, -749, -7938, 29843, 11073, 5531}, '{26611, -6428, 17315, -22263, 13033, -24563, -11851, 23878, -19496}, '{25354, -12167, -31445, -4507, 30085, 20648, -31500, -11505, 25614}, '{-22059, -8192, -10973, -10655, -12914, 18182, 25176, 11766, -11261}, '{-31420, 1125, 15848, 23391, 18331, -28046, -6167, 23107, 7970}, '{8617, 4877, 8063, 9329, -5743, -16022, -9560, -25107, -7222}, '{-25818, 15914, 4419, 13595, 28604, -11633, -17678, 30626, 7652}, '{17130, -409, 3762, 6188, -7852, -32204, 18329, 32459, 4268}, '{-28591, 32767, -7547, 30291, -32057, 28927, 5956, 24159, 27997}},
        '{'{-32662, 754, 1627, -2912, -25109, 937, -21294, 4509, -115}, '{4082, -27284, -5495, -12234, 27528, 23577, -5983, -24047, 12785}, '{18863, 28176, 13873, -29634, -19641, 24414, 20478, -9264, 9302}, '{-22021, 22693, -15095, 12206, -28020, 13400, -2691, -31371, -5738}, '{-840, 15950, -5587, -30943, -15682, -9724, -13499, -28035, 5196}, '{681, 10636, 24320, 11973, 30870, -30999, 23905, 19121, -397}, '{28481, 10634, -20282, 30842, 30736, 15047, -9829, 23846, -14229}, '{31828, 30121, -19758, -28045, 24554, -28218, -29786, 32418, 6257}, '{-3382, -4353, 20839, -22744, 40, -101, -12194, -4101, 23716}},
        '{'{-6046, 12859, 27225, 1947, 696, -25473, -3142, -31457, -29904}, '{-25621, 26750, 4483, 28992, -475, 20983, -14681, -11252, -21676}, '{3531, -18100, 5752, -28302, -37, -11345, 4409, 18581, 28524}, '{524, 22511, 17041, -9817, -24673, -22929, -26979, 6583, 2497}, '{9509, -17920, -23785, -27763, 136, -17964, -18379, -30510, 31056}, '{12045, -18040, 11654, -7781, -21339, 419, -472, 28314, 6494}, '{-31796, -583, -14035, -28848, -4806, 7319, -13570, 23794, -32022}, '{-31800, 8183, -1034, -13872, -4875, 11133, -18926, -27702, -30833}, '{25062, -26755, -27816, -2076, 22255, 19264, -25213, 20442, 19348}}
    },
    '{
        '{'{5103, 11439, 18878, 29025, 3096, 27346, -2264, -18295, -19128}, '{27847, 32220, 6127, 16681, -2285, -9514, 9539, 30711, -26674}, '{11391, 28279, 8002, -18729, -12053, -27624, -12716, -10589, 30586}, '{19886, 4640, -19678, 22058, 860, 6181, 16612, -3246, -15305}, '{-26774, -21981, -16409, 16739, 23617, 14685, 13972, -27419, 18787}, '{-19666, 7522, 91, 30782, 26686, -24079, 18683, -21938, 4970}, '{-18274, -17061, -20429, -9724, 14020, 902, 16105, -215, 7427}, '{2727, -22036, 23652, 6555, 16013, 16684, 6400, -22710, -29987}, '{-31922, -31616, -13056, -26528, 18292, -16629, -10211, 23941, 18501}},
        '{'{-11591, -23266, -5358, 4714, -8176, -6281, 11601, 13515, -22519}, '{-14455, -9510, -7092, 26304, -27417, -6244, -14602, 11085, 29527}, '{11194, 10873, 7600, -4709, -22677, -3943, -26668, -10129, -10676}, '{-14824, -12539, -19422, -16308, 11451, -29141, 9167, -23749, 3349}, '{7652, -25103, 6654, -26260, -14836, -21648, 31842, 25221, 16148}, '{-31108, -1377, 30562, 26903, -2541, -26027, -29905, -30726, 20230}, '{68, -11063, 32280, 13231, -8288, 6090, 27354, -11813, 1296}, '{-31006, -9066, -27523, -15332, -20196, 2673, 24526, -25755, -21927}, '{-15227, 17986, -10845, 25291, 15283, 19021, -10269, 27320, -8737}},
        '{'{21982, 23813, 26653, 22619, 30713, -16459, 29121, -2755, 20968}, '{19610, -25316, 999, -13913, 15969, 105, 23215, -18323, -2144}, '{20857, -20220, 21942, 2432, -7925, 8371, 16995, -15420, -8422}, '{-497, -9743, -7460, 31594, 21392, 29556, -7098, -5384, 26719}, '{17410, 12796, 32017, -21262, 12097, 14496, -30495, 9638, 2628}, '{-14498, -25340, -3077, -14001, 21631, 20757, -28807, 30067, 9318}, '{30474, -20208, -30718, 14126, 17085, 22702, 21614, -14048, 24807}, '{-18537, -28995, -7807, -21212, 3929, 264, 22063, 27483, 17408}, '{-32605, 23578, -27458, -26769, 2996, -16406, 9878, 23199, 3713}}
    },
    '{
        '{'{-6307, 2307, -32509, 9570, -27532, 24740, 22954, -3730, 13332}, '{-27415, -14203, 31448, 25599, -5037, 25270, 13029, 19715, -4269}, '{29847, 27696, -17570, -15714, -15143, -18553, 16298, -15732, 7684}, '{-20240, -19557, 4300, -16785, -11574, 32508, 16811, -4427, 4334}, '{28298, 2803, -8149, 26374, 711, 14848, -7629, -15710, 31584}, '{31767, 13760, 30407, -98, 8978, 13088, -16382, -8538, -29428}, '{-31168, 4990, 17148, 27720, -14589, -17011, -3202, 2010, -28541}, '{9446, 27078, 20102, 22932, 4922, 26626, 981, 24751, 9727}, '{-29004, -29126, -12178, -10670, 12542, -2480, -22215, 16043, -2783}},
        '{'{-25110, -12219, -4899, 13391, 7257, -15891, -21515, -27368, 4452}, '{-21828, -31879, 27456, -2627, 21581, -23028, -19770, 1137, -13775}, '{8323, 21408, -29581, -31055, 20195, 27021, -32693, -13295, 16452}, '{-4649, -26321, -32438, 22950, -25996, -13067, -15514, -18000, -14812}, '{5597, 29465, 8739, -29241, -15424, -18624, 1032, 3011, -5370}, '{-5019, -29700, -29305, 29619, -25139, 82, 10616, -6639, -28925}, '{11390, 7432, -8145, -18901, 11965, -14589, 20780, -14261, 16373}, '{22833, -23502, -17270, 25771, -11569, -3109, 3174, -28098, 7651}, '{22866, 28413, 19774, -14987, -13917, -20139, 924, -11333, -26399}},
        '{'{-11175, -32310, -14847, -3590, -25195, 21401, 20106, -13704, 17833}, '{-3059, -4429, -4798, 18642, 5332, -14713, -21720, -24264, -7851}, '{14373, 5550, -11053, -23078, 9911, -29306, 15872, 17800, 7164}, '{23253, 15739, -12049, 17061, 21443, 686, -15640, -15959, 17244}, '{-29633, 5177, 25591, -24988, 6695, 4801, 9651, 17085, 29037}, '{-10555, -23622, -165, 8543, 17320, 30793, -13643, 32632, 2567}, '{-24221, 27567, -7483, 25257, -23780, -8970, -9350, 19285, -27893}, '{4611, -14062, 6051, 24622, -18071, -17263, -7057, 22683, -23498}, '{23151, -19767, -13933, 28871, -8633, -4251, -4693, 22526, -15444}}
    },
    '{
        '{'{9838, -20818, -30046, -3423, -1974, -28297, 11077, -17956, 26414}, '{-23648, 4307, 17831, 20894, -13089, 1903, -19281, -20607, -4192}, '{-19586, 1128, 22897, -23873, 21623, 7469, 2231, -19346, -8330}, '{11584, 869, -29227, -8554, -27237, 26629, 24429, 1059, -27795}, '{7971, 30332, 21096, -9021, 19612, -20901, -24837, -6007, 16683}, '{9859, -20373, 3979, 32691, -6698, -5526, 1770, -8060, 26269}, '{-16068, 6572, 24578, -21538, 17477, 9775, -23348, 18065, 2127}, '{-5448, 13865, 21400, 15061, -24984, -23037, 3772, 16174, 18800}, '{1183, 12742, -22529, -24781, 97, -21329, 11531, -14489, -23234}},
        '{'{-24952, 10430, 7299, 13239, -26517, -2250, 10983, -8023, -10954}, '{-12007, 20333, 10630, -16313, 3816, -7233, 21853, -23810, 20421}, '{-23002, -30781, -31481, 16754, -85, -27753, -29480, -12302, 29469}, '{-10957, 16273, 9912, -6869, -25695, -1232, -21810, 2922, -3670}, '{-24880, -28433, 14325, 11393, -662, 6709, 13760, 27379, 25983}, '{25656, 21647, -32432, 12488, -11927, 9876, 14013, 12479, -17610}, '{1451, -28263, 128, -26501, 31025, 2471, -32382, -15162, 19331}, '{-4322, -23795, 30484, 884, -8885, 32011, -17787, 8048, -32112}, '{14797, -15170, -8824, -24549, -27770, -1684, 28406, -11734, -13692}},
        '{'{-9240, 3817, -24177, 18364, 15744, -17241, -8667, 4614, -20749}, '{29277, 19258, 30575, -30823, -31156, 30784, 29630, -16460, -28622}, '{16561, -31332, 9210, -17465, -13887, 3692, 28400, -7118, -13945}, '{26600, -20710, 32424, 10557, 2736, -11794, -15210, 782, -7873}, '{13791, 1877, 21044, 16775, 3108, 28112, -8506, -21270, 2452}, '{18982, -9852, 30864, -6430, -17297, 27832, 16635, 29551, 25358}, '{13295, 21223, -21377, -26609, -8744, 8846, -26742, -27914, 7428}, '{-19884, 29801, -17688, 564, 11979, 11516, 20277, 26077, -31933}, '{10484, -6356, -23334, 19836, -20261, -22782, 2236, -6078, -13827}}
    },
    '{
        '{'{23063, -19731, 6172, -1799, 31541, 15250, 14191, -4165, 3649}, '{17476, 5156, -2223, -23528, 31449, -20629, 11596, 12578, -25259}, '{31544, 22514, -8641, 26569, 17700, 24427, 22953, 12550, 19345}, '{-9953, -7686, -6542, 30959, 5100, 15878, 178, 8976, 16158}, '{7964, -13185, -24117, 160, 10086, 20953, 21030, -18147, 32002}, '{-2477, -7860, -6254, 25664, 27049, -15210, 31249, 12970, 10244}, '{-26492, 17810, 10949, 26638, -32758, 24882, 5085, -29997, 11042}, '{16387, 7176, -25638, 1618, -8636, 27271, -26262, -25251, -29661}, '{-16689, -3026, -851, -17981, -28102, -11645, 18630, -25534, 11237}},
        '{'{-19816, 1719, -9797, -26973, -11005, 32327, -101, -29710, 19266}, '{5630, -18064, -15801, 3082, -6035, -27457, -25221, 10352, 21881}, '{-24571, -16908, -25304, -42, 8628, -2133, 19905, 13190, -16612}, '{-32379, 24808, 1610, 29319, -6371, -1180, 24914, -4049, -30276}, '{-26305, -25989, 31170, -24279, 22045, -19360, 28209, -13636, -11468}, '{21017, -476, -15725, -24736, -6923, -7589, -13158, -25032, 23864}, '{-28900, -16467, -29737, 8658, 32005, 17345, -26027, -13022, 13185}, '{-23971, 22253, 18402, 14606, -3862, -6626, 26505, -5706, -28901}, '{-32377, 24524, -25251, 20132, 20646, -24484, 15985, -18859, -26409}},
        '{'{-6747, 3988, 781, -12179, 9896, -590, -29207, -1738, -21378}, '{-2623, -17592, 4154, -22425, 29548, -23479, -13775, 4369, -7887}, '{-23463, -17961, 3001, 11240, -20231, -3981, 4810, -13478, -8947}, '{26911, 11388, 32277, -27807, 18925, 6401, 21984, -1877, -5449}, '{838, 3362, -19490, 23086, 22874, 9702, 31716, -7535, -1168}, '{5388, 15924, 31535, -23180, 9127, 6000, 31664, -28745, -9575}, '{31552, 8508, 17382, -19298, 10473, -2321, -9116, 24166, -17572}, '{31210, 7895, -9649, 29094, -666, 12246, 16176, -27385, 27173}, '{-1806, -10430, 30797, 1300, 11054, -24099, -32480, -18636, 10679}}
    }
};
