logic signed [7:0] convolve11_weight[4][8][3][3] = '{
    '{
        '{'{92, -81, -80}, '{-9, 71, -11}, '{-61, -5, 71}},
        '{'{-66, 72, -91}, '{-123, -31, -73}, '{92, 46, -90}},
        '{'{-79, -120, -6}, '{65, -62, -66}, '{-112, 61, 66}},
        '{'{-117, 31, 10}, '{-108, -28, -114}, '{-8, -76, 71}},
        '{'{29, 5, -114}, '{-14, 110, 79}, '{-77, -96, 23}},
        '{'{121, -37, -122}, '{73, -8, -63}, '{-53, -41, 124}},
        '{'{70, -88, 60}, '{-92, 12, 35}, '{-66, 69, -66}},
        '{'{58, -52, -110}, '{0, -127, 84}, '{77, -38, -16}}
    },
    '{
        '{'{-21, 21, -50}, '{-115, 104, -61}, '{-23, 17, -123}},
        '{'{-102, 63, 27}, '{107, 109, 41}, '{-115, -83, 48}},
        '{'{-72, -70, -111}, '{86, -33, 89}, '{92, 77, 7}},
        '{'{-102, -111, 68}, '{-85, 47, 94}, '{-3, -36, 121}},
        '{'{-56, 58, -101}, '{-122, 7, 53}, '{-9, 120, -102}},
        '{'{-5, 75, -91}, '{-35, 49, -108}, '{93, -9, 56}},
        '{'{61, 55, 92}, '{23, 57, 9}, '{0, -26, 19}},
        '{'{71, -78, -90}, '{67, 124, 30}, '{-91, 56, -2}}
    },
    '{
        '{'{105, 5, -69}, '{80, 90, 61}, '{-97, 70, -39}},
        '{'{75, 17, -97}, '{31, -44, -38}, '{-89, 117, 50}},
        '{'{-54, -90, -60}, '{-5, -89, -1}, '{79, -115, 35}},
        '{'{102, -5, 11}, '{-25, -53, 112}, '{-74, 36, -46}},
        '{'{75, 51, 34}, '{58, -48, -100}, '{9, -27, -120}},
        '{'{17, 112, 108}, '{92, 25, -34}, '{-5, -27, 59}},
        '{'{-5, 94, 121}, '{-69, 58, -110}, '{-116, 1, -101}},
        '{'{-118, 67, 61}, '{-112, -101, -4}, '{-122, -128, -121}}
    },
    '{
        '{'{25, -61, -69}, '{120, -12, 127}, '{36, 44, 85}},
        '{'{-15, 118, 127}, '{72, -17, 38}, '{42, 97, 36}},
        '{'{-60, -37, -115}, '{13, 41, -56}, '{6, -34, 12}},
        '{'{-30, 3, 104}, '{-112, -123, -88}, '{55, 29, 53}},
        '{'{-106, -27, -105}, '{123, -6, 36}, '{107, 59, -94}},
        '{'{70, 6, -40}, '{-52, -111, -33}, '{-80, -91, -128}},
        '{'{74, -15, -20}, '{-124, -33, 60}, '{-1, -118, -99}},
        '{'{-31, -23, 112}, '{-115, -109, -87}, '{76, 44, -77}}
    }
};
