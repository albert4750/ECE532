localparam bit signed [0:2][0:26][19:0] Input1 = '{
    '{-20'd97, -20'd8, -20'd127, -20'd63, 20'd103, 20'd41, -20'd71, -20'd93, -20'd26, -20'd9, -20'd117, 20'd46, -20'd46, -20'd37, 20'd0, 20'd14, -20'd29, -20'd75, 20'd12, -20'd7, 20'd42, -20'd44, 20'd75, -20'd60, -20'd122, 20'd68, -20'd81},
    '{-20'd1, 20'd116, 20'd3, 20'd76, -20'd28, 20'd52, 20'd104, -20'd50, 20'd15, 20'd20, 20'd99, 20'd58, -20'd105, 20'd79, 20'd13, -20'd11, -20'd43, -20'd80, -20'd79, -20'd59, 20'd41, 20'd35, 20'd64, -20'd33, 20'd69, -20'd34, -20'd128},
    '{-20'd15, 20'd50, -20'd92, 20'd34, -20'd80, -20'd35, 20'd3, -20'd30, -20'd86, 20'd77, -20'd16, 20'd103, 20'd21, 20'd73, -20'd1, -20'd128, 20'd10, -20'd14, -20'd85, 20'd58, -20'd1, -20'd105, 20'd59, 20'd2, -20'd7, -20'd30, -20'd66}
};
