localparam bit signed [0:2][0:31][0:4][0:4][24:0] Weight3 = '{
    '{'{'{25'd42540, 25'd9116, 25'd1519, 25'd16712, 25'd15193}, '{25'd47098, -25'd1519, 25'd25828, 25'd9116, 25'd9116}, '{25'd41021, 25'd9116, 25'd13674, 25'd3039, 25'd22789}, '{25'd31905, 25'd12154, 25'd18232, -25'd7596, 25'd25828}, '{25'd57733, 25'd3039, 25'd13674, 25'd10635, 25'd21270}}, '{'{25'd6077, 25'd25828, 25'd18232, 25'd27347, 25'd25828}, '{25'd22789, 25'd3039, 25'd9116, -25'd3039, 25'd10635}, '{25'd9116, -25'd3039, 25'd10635, -25'd3039, 25'd34944}, '{25'd24309, 25'd13674, 25'd19751, 25'd22789, 25'd37982}, '{25'd44060, 25'd37982, 25'd31905, 25'd53175, 25'd69888}}, '{'{25'd112428, 25'd63811, 25'd59253, 25'd60772, 25'd95716}, '{25'd62291, 25'd25828, 25'd28867, 25'd12154, 25'd53175}, '{25'd69888, 25'd16712, 25'd44060, 25'd37982, 25'd65330}, '{25'd47098, 25'd13674, 25'd16712, 25'd10635, 25'd59253}, '{25'd57733, 25'd34944, 25'd34944, 25'd34944, 25'd60772}}, '{'{-25'd53175, -25'd30386, -25'd42540, -25'd19751, -25'd36463}, '{-25'd54695, -25'd37982, -25'd25828, -25'd33425, -25'd36463}, '{-25'd53175, -25'd24309, -25'd10635, -25'd34944, -25'd37982}, '{-25'd53175, -25'd31905, -25'd16712, -25'd13674, -25'd28867}, '{-25'd80523, -25'd54695, -25'd36463, -25'd56214, -25'd59253}}, '{'{25'd21270, 25'd22789, 25'd25828, 25'd24309, 25'd37982}, '{25'd16712, 25'd12154, 25'd19751, 25'd16712, 25'd19751}, '{25'd33425, 25'd21270, 25'd18232, 25'd28867, 25'd16712}, '{25'd33425, 25'd10635, 25'd15193, 25'd18232, 25'd31905}, '{25'd56214, 25'd31905, 25'd57733, 25'd45579, 25'd89639}}, '{'{25'd25828, 25'd30386, 25'd16712, 25'd24309, 25'd45579}, '{25'd37982, 25'd28867, 25'd28867, 25'd15193, 25'd31905}, '{25'd34944, 25'd10635, 25'd0, 25'd18232, 25'd30386}, '{25'd9116, 25'd1519, 25'd3039, 25'd0, 25'd19751}, '{25'd1519, 25'd3039, -25'd4558, -25'd9116, 25'd3039}}, '{'{-25'd9116, -25'd34944, -25'd13674, -25'd15193, 25'd1519}, '{-25'd9116, -25'd31905, -25'd16712, -25'd13674, -25'd10635}, '{-25'd10635, -25'd33425, -25'd12154, -25'd18232, -25'd15193}, '{-25'd30386, -25'd19751, -25'd10635, -25'd27347, -25'd12154}, '{25'd6077, -25'd13674, -25'd18232, -25'd21270, 25'd4558}}, '{'{25'd6077, -25'd10635, -25'd15193, -25'd18232, -25'd18232}, '{-25'd16712, 25'd6077, -25'd19751, 25'd0, -25'd12154}, '{-25'd9116, -25'd31905, -25'd19751, -25'd27347, -25'd33425}, '{-25'd30386, -25'd19751, -25'd36463, -25'd37982, -25'd36463}, '{-25'd27347, -25'd50137, -25'd25828, -25'd45579, -25'd37982}}, '{'{25'd91158, 25'd48618, 25'd50137, 25'd51656, 25'd92677}, '{25'd72926, 25'd10635, 25'd31905, 25'd22789, 25'd68368}, '{25'd74446, 25'd37982, 25'd13674, 25'd28867, 25'd75965}, '{25'd68368, 25'd41021, 25'd27347, 25'd27347, 25'd83561}, '{25'd98754, 25'd48618, 25'd48618, 25'd63811, 25'd106351}}, '{'{-25'd24309, -25'd1519, 25'd16712, 25'd7596, 25'd16712}, '{-25'd12154, 25'd1519, 25'd33425, 25'd28867, 25'd24309}, '{25'd13674, 25'd21270, 25'd10635, 25'd12154, 25'd6077}, '{25'd9116, 25'd18232, 25'd33425, 25'd18232, 25'd18232}, '{25'd12154, 25'd25828, 25'd36463, 25'd7596, 25'd24309}}, '{'{25'd91158, 25'd27347, 25'd25828, 25'd39502, 25'd68368}, '{25'd50137, 25'd15193, -25'd4558, 25'd12154, 25'd31905}, '{25'd48618, 25'd6077, 25'd7596, -25'd3039, 25'd27347}, '{25'd54695, 25'd6077, -25'd22789, -25'd7596, 25'd34944}, '{25'd120025, 25'd54695, 25'd37982, 25'd36463, 25'd94197}}, '{'{-25'd60772, -25'd53175, -25'd39502, -25'd56214, -25'd54695}, '{-25'd37982, -25'd31905, -25'd15193, -25'd22789, -25'd41021}, '{-25'd36463, -25'd25828, -25'd27347, -25'd33425, -25'd37982}, '{-25'd42540, -25'd16712, -25'd31905, -25'd34944, -25'd48618}, '{-25'd59253, -25'd24309, -25'd16712, -25'd42540, -25'd48618}}, '{'{25'd0, 25'd0, 25'd24309, 25'd4558, -25'd22789}, '{25'd10635, 25'd22789, 25'd19751, 25'd0, -25'd4558}, '{-25'd4558, 25'd25828, 25'd28867, 25'd6077, 25'd4558}, '{25'd9116, 25'd10635, 25'd7596, 25'd31905, 25'd1519}, '{-25'd4558, 25'd16712, 25'd22789, 25'd1519, -25'd7596}}, '{'{-25'd36463, -25'd16712, -25'd1519, -25'd10635, 25'd0}, '{-25'd21270, -25'd10635, -25'd22789, -25'd16712, -25'd12154}, '{-25'd9116, 25'd0, -25'd9116, 25'd1519, -25'd19751}, '{-25'd12154, -25'd13674, -25'd10635, -25'd3039, -25'd18232}, '{25'd1519, 25'd0, 25'd1519, 25'd0, -25'd3039}}, '{'{25'd34944, 25'd25828, 25'd31905, 25'd16712, 25'd39502}, '{25'd18232, 25'd4558, 25'd21270, 25'd12154, 25'd41021}, '{25'd36463, 25'd28867, 25'd25828, 25'd30386, 25'd30386}, '{25'd19751, 25'd19751, 25'd4558, 25'd6077, 25'd34944}, '{25'd37982, 25'd41021, 25'd28867, 25'd53175, 25'd62291}}, '{'{25'd4558, 25'd6077, 25'd25828, 25'd9116, 25'd37982}, '{25'd27347, -25'd1519, 25'd1519, 25'd27347, 25'd27347}, '{25'd12154, 25'd24309, 25'd4558, 25'd33425, 25'd28867}, '{25'd25828, 25'd24309, 25'd34944, 25'd18232, 25'd31905}, '{25'd42540, 25'd42540, 25'd41021, 25'd57733, 25'd56214}}, '{'{25'd135218, 25'd88119, 25'd98754, 25'd100274, 25'd121544}, '{25'd85081, 25'd45579, 25'd71407, 25'd50137, 25'd80523}, '{25'd80523, 25'd57733, 25'd56214, 25'd54695, 25'd74446}, '{25'd85081, 25'd48618, 25'd72926, 25'd65330, 25'd65330}, '{25'd123063, 25'd91158, 25'd89639, 25'd80523, 25'd85081}}, '{'{-25'd3039, -25'd22789, -25'd28867, -25'd47098, -25'd88119}, '{-25'd22789, -25'd18232, -25'd10635, -25'd22789, -25'd28867}, '{-25'd1519, -25'd21270, -25'd9116, -25'd1519, -25'd28867}, '{-25'd28867, -25'd24309, -25'd12154, -25'd24309, -25'd7596}, '{-25'd16712, -25'd16712, -25'd9116, -25'd18232, -25'd19751}}, '{'{-25'd51656, -25'd15193, -25'd7596, -25'd37982, -25'd62291}, '{-25'd31905, -25'd15193, -25'd19751, -25'd15193, -25'd47098}, '{-25'd45579, -25'd3039, 25'd15193, -25'd7596, -25'd27347}, '{-25'd44060, -25'd22789, 25'd10635, -25'd16712, -25'd41021}, '{-25'd72926, -25'd31905, -25'd30386, -25'd18232, -25'd62291}}, '{'{25'd92677, 25'd54695, 25'd71407, 25'd65330, 25'd97235}, '{25'd82042, 25'd28867, 25'd30386, 25'd51656, 25'd68368}, '{25'd57733, 25'd33425, 25'd16712, 25'd31905, 25'd63811}, '{25'd79004, 25'd34944, 25'd45579, 25'd37982, 25'd66849}, '{25'd101793, 25'd85081, 25'd74446, 25'd72926, 25'd109390}}, '{'{-25'd50137, -25'd37982, -25'd34944, -25'd30386, -25'd37982}, '{-25'd53175, -25'd34944, -25'd15193, -25'd16712, -25'd41021}, '{-25'd41021, -25'd25828, -25'd30386, -25'd34944, -25'd47098}, '{-25'd51656, -25'd30386, -25'd41021, -25'd21270, -25'd47098}, '{-25'd59253, -25'd34944, -25'd25828, -25'd39502, -25'd42540}}, '{'{25'd189912, 25'd144333, 25'd150411, 25'd158007, 25'd191432}, '{25'd145853, 25'd113947, 25'd101793, 25'd115467, 25'd139776}, '{25'd156488, 25'd92677, 25'd95716, 25'd103312, 25'd138256}, '{25'd144333, 25'd116986, 25'd100274, 25'd83561, 25'd138256}, '{25'd192951, 25'd144333, 25'd135218, 25'd116986, 25'd148891}}, '{'{-25'd113947, -25'd75965, -25'd60772, -25'd57733, -25'd74446}, '{-25'd47098, -25'd22789, 25'd0, -25'd18232, -25'd57733}, '{-25'd41021, -25'd16712, -25'd15193, 25'd3039, -25'd28867}, '{-25'd27347, -25'd15193, -25'd16712, -25'd30386, -25'd60772}, '{-25'd9116, -25'd15193, 25'd1519, -25'd6077, -25'd41021}}, '{'{25'd12154, 25'd21270, 25'd27347, 25'd4558, 25'd27347}, '{-25'd15193, -25'd1519, -25'd15193, -25'd7596, -25'd4558}, '{-25'd18232, 25'd1519, -25'd15193, -25'd1519, 25'd0}, '{-25'd6077, 25'd7596, -25'd7596, -25'd4558, 25'd10635}, '{25'd10635, 25'd6077, -25'd9116, 25'd10635, 25'd3039}}, '{'{25'd44060, 25'd30386, 25'd33425, 25'd48618, 25'd91158}, '{25'd19751, 25'd31905, 25'd25828, 25'd25828, 25'd54695}, '{25'd24309, 25'd15193, 25'd9116, 25'd31905, 25'd50137}, '{25'd45579, 25'd22789, 25'd15193, 25'd45579, 25'd63811}, '{25'd74446, 25'd54695, 25'd62291, 25'd85081, 25'd118505}}, '{'{25'd33425, 25'd18232, 25'd16712, 25'd3039, 25'd28867}, '{25'd16712, 25'd7596, 25'd16712, 25'd7596, 25'd30386}, '{25'd19751, 25'd22789, 25'd21270, 25'd9116, 25'd39502}, '{25'd15193, 25'd9116, 25'd16712, 25'd13674, 25'd27347}, '{25'd15193, 25'd30386, 25'd30386, 25'd22789, 25'd33425}}, '{'{25'd75965, 25'd37982, 25'd28867, 25'd44060, 25'd66849}, '{25'd50137, 25'd51656, 25'd30386, 25'd37982, 25'd34944}, '{25'd48618, 25'd33425, 25'd44060, 25'd44060, 25'd57733}, '{25'd66849, 25'd51656, 25'd37982, 25'd31905, 25'd33425}, '{25'd36463, 25'd13674, 25'd13674, 25'd16712, 25'd33425}}, '{'{25'd10635, -25'd7596, 25'd3039, 25'd4558, 25'd31905}, '{25'd4558, -25'd19751, -25'd24309, -25'd18232, 25'd22789}, '{25'd21270, -25'd19751, -25'd27347, -25'd24309, 25'd15193}, '{25'd10635, -25'd12154, -25'd9116, -25'd22789, 25'd15193}, '{25'd65330, 25'd13674, 25'd36463, 25'd36463, 25'd72926}}, '{'{25'd95716, 25'd54695, 25'd60772, 25'd62291, 25'd100274}, '{25'd72926, 25'd19751, 25'd28867, 25'd24309, 25'd79004}, '{25'd71407, 25'd16712, 25'd30386, 25'd24309, 25'd68368}, '{25'd94197, 25'd51656, 25'd30386, 25'd34944, 25'd75965}, '{25'd98754, 25'd82042, 25'd63811, 25'd51656, 25'd100274}}, '{'{25'd39502, 25'd25828, 25'd4558, 25'd3039, 25'd48618}, '{25'd37982, -25'd3039, 25'd3039, 25'd18232, 25'd21270}, '{25'd28867, 25'd16712, 25'd1519, 25'd1519, 25'd36463}, '{25'd18232, 25'd4558, 25'd7596, 25'd1519, 25'd28867}, '{25'd28867, 25'd10635, 25'd9116, 25'd9116, 25'd42540}}, '{'{25'd150411, 25'd72926, 25'd69888, 25'd71407, 25'd145853}, '{25'd95716, 25'd24309, 25'd21270, 25'd25828, 25'd92677}, '{25'd66849, 25'd3039, -25'd1519, 25'd22789, 25'd65330}, '{25'd86600, 25'd31905, 25'd1519, 25'd16712, 25'd88119}, '{25'd138256, 25'd91158, 25'd59253, 25'd75965, 25'd167123}}, '{'{25'd59253, 25'd6077, 25'd15193, 25'd24309, 25'd28867}, '{25'd59253, 25'd3039, -25'd7596, 25'd16712, 25'd27347}, '{25'd34944, 25'd13674, 25'd4558, 25'd10635, 25'd13674}, '{25'd50137, 25'd16712, 25'd18232, 25'd6077, 25'd13674}, '{25'd63811, 25'd13674, 25'd39502, 25'd36463, 25'd22789}}},
    '{'{'{25'd9728, 25'd9728, 25'd9728, 25'd0, 25'd32428}, '{-25'd3243, 25'd8107, 25'd8107, -25'd4864, 25'd14592}, '{-25'd1621, 25'd14592, 25'd1621, 25'd0, 25'd21078}, '{25'd4864, 25'd1621, -25'd3243, 25'd1621, 25'd19457}, '{25'd6486, 25'd1621, 25'd11350, 25'd25942, 25'd25942}}, '{'{25'd21078, 25'd37292, 25'd3243, 25'd19457, 25'd19457}, '{25'd34049, 25'd27564, -25'd4864, 25'd29185, 25'd11350}, '{25'd24321, 25'd11350, -25'd8107, 25'd11350, -25'd1621}, '{25'd16214, 25'd17835, 25'd0, 25'd16214, 25'd16214}, '{-25'd14592, -25'd6486, -25'd3243, -25'd14592, 25'd9728}}, '{'{-25'd56749, -25'd43777, -25'd42156, -25'd38913, -25'd53506}, '{-25'd50263, -25'd17835, -25'd16214, -25'd37292, -25'd37292}, '{-25'd29185, -25'd12971, -25'd21078, -25'd21078, -25'd38913}, '{-25'd32428, -25'd27564, -25'd32428, -25'd16214, -25'd30806}, '{-25'd68098, -25'd45399, -25'd35671, -25'd48642, -25'd51884}}, '{'{25'd69720, 25'd59991, 25'd50263, 25'd48642, 25'd43777}, '{25'd53506, 25'd37292, 25'd35671, 25'd21078, 25'd42156}, '{25'd69720, 25'd27564, 25'd29185, 25'd16214, 25'd42156}, '{25'd63234, 25'd35671, 25'd14592, 25'd43777, 25'd55127}, '{25'd84312, 25'd63234, 25'd50263, 25'd58370, 25'd72962}}, '{'{-25'd9728, -25'd29185, -25'd32428, -25'd21078, -25'd40535}, '{-25'd16214, 25'd1621, -25'd24321, -25'd19457, -25'd43777}, '{-25'd9728, -25'd16214, -25'd19457, -25'd8107, -25'd42156}, '{-25'd14592, -25'd19457, -25'd34049, -25'd35671, -25'd47020}, '{-25'd56749, -25'd64856, -25'd43777, -25'd53506, -25'd79448}}, '{'{-25'd14592, 25'd4864, -25'd16214, -25'd4864, 25'd8107}, '{-25'd21078, -25'd9728, 25'd4864, 25'd1621, -25'd9728}, '{25'd4864, -25'd9728, -25'd6486, -25'd4864, 25'd9728}, '{-25'd16214, -25'd8107, 25'd6486, -25'd6486, -25'd4864}, '{25'd6486, 25'd4864, 25'd9728, 25'd1621, 25'd32428}}, '{'{25'd32428, 25'd43777, 25'd22699, 25'd12971, 25'd19457}, '{25'd25942, 25'd32428, 25'd17835, 25'd11350, 25'd25942}, '{25'd22699, 25'd30806, 25'd29185, 25'd8107, 25'd17835}, '{25'd27564, 25'd24321, 25'd27564, 25'd24321, 25'd21078}, '{25'd45399, 25'd48642, 25'd29185, 25'd17835, 25'd11350}}, '{'{25'd50263, 25'd34049, 25'd24321, 25'd25942, 25'd55127}, '{25'd24321, 25'd29185, 25'd1621, 25'd21078, 25'd35671}, '{25'd32428, 25'd27564, 25'd12971, 25'd29185, 25'd40535}, '{25'd45399, 25'd27564, 25'd29185, 25'd35671, 25'd42156}, '{25'd77827, 25'd47020, 25'd58370, 25'd58370, 25'd71341}}, '{'{-25'd79448, -25'd29185, -25'd38913, -25'd50263, -25'd77827}, '{-25'd64856, -25'd29185, -25'd9728, -25'd11350, -25'd51884}, '{-25'd40535, -25'd22699, -25'd6486, -25'd32428, -25'd55127}, '{-25'd68098, -25'd25942, -25'd22699, -25'd17835, -25'd56749}, '{-25'd69720, -25'd56749, -25'd30806, -25'd47020, -25'd81069}}, '{'{25'd3243, -25'd16214, -25'd21078, -25'd16214, -25'd4864}, '{-25'd4864, -25'd17835, -25'd19457, -25'd21078, -25'd37292}, '{-25'd24321, -25'd27564, -25'd32428, -25'd27564, -25'd25942}, '{-25'd17835, -25'd9728, -25'd30806, -25'd6486, -25'd14592}, '{-25'd4864, -25'd22699, -25'd29185, -25'd17835, -25'd19457}}, '{'{-25'd110254, -25'd59991, -25'd63234, -25'd53506, -25'd81069}, '{-25'd64856, -25'd48642, -25'd34049, -25'd30806, -25'd71341}, '{-25'd69720, -25'd35671, -25'd22699, -25'd45399, -25'd50263}, '{-25'd43777, -25'd30806, -25'd14592, -25'd17835, -25'd40535}, '{-25'd105390, -25'd63234, -25'd64856, -25'd56749, -25'd81069}}, '{'{25'd97283, 25'd59991, 25'd50263, 25'd59991, 25'd116740}, '{25'd51884, 25'd27564, 25'd8107, 25'd8107, 25'd64856}, '{25'd63234, 25'd38913, 25'd8107, 25'd37292, 25'd53506}, '{25'd37292, 25'd29185, 25'd16214, 25'd11350, 25'd64856}, '{25'd69720, 25'd42156, 25'd37292, 25'd34049, 25'd76205}}, '{'{25'd50263, 25'd6486, 25'd22699, 25'd9728, 25'd69720}, '{25'd8107, 25'd9728, -25'd6486, -25'd11350, 25'd17835}, '{25'd12971, 25'd4864, -25'd8107, 25'd6486, 25'd12971}, '{25'd34049, -25'd14592, -25'd21078, -25'd3243, 25'd17835}, '{25'd34049, 25'd29185, 25'd24321, 25'd16214, 25'd58370}}, '{'{25'd19457, 25'd8107, 25'd25942, 25'd24321, 25'd29185}, '{25'd27564, 25'd12971, -25'd6486, 25'd14592, 25'd3243}, '{25'd30806, 25'd24321, 25'd17835, 25'd6486, 25'd22699}, '{25'd32428, 25'd0, -25'd6486, -25'd8107, 25'd21078}, '{25'd14592, 25'd16214, -25'd8107, 25'd8107, -25'd6486}}, '{'{-25'd51884, -25'd43777, -25'd40535, -25'd38913, -25'd81069}, '{-25'd58370, -25'd25942, -25'd16214, -25'd30806, -25'd40535}, '{-25'd29185, -25'd14592, -25'd22699, -25'd22699, -25'd37292}, '{-25'd56749, -25'd12971, -25'd22699, -25'd11350, -25'd47020}, '{-25'd50263, -25'd29185, -25'd42156, -25'd34049, -25'd69720}}, '{'{-25'd22699, -25'd11350, -25'd3243, -25'd25942, -25'd25942}, '{-25'd3243, -25'd9728, -25'd17835, -25'd17835, -25'd32428}, '{-25'd22699, -25'd16214, -25'd21078, -25'd19457, -25'd34049}, '{-25'd16214, -25'd12971, -25'd11350, -25'd30806, -25'd30806}, '{-25'd40535, -25'd34049, -25'd40535, -25'd25942, -25'd47020}}, '{'{-25'd84312, -25'd50263, -25'd63234, -25'd50263, -25'd69720}, '{-25'd48642, -25'd34049, -25'd48642, -25'd47020, -25'd42156}, '{-25'd51884, -25'd40535, -25'd30806, -25'd21078, -25'd32428}, '{-25'd47020, -25'd40535, -25'd24321, -25'd22699, -25'd59991}, '{-25'd81069, -25'd50263, -25'd51884, -25'd55127, -25'd71341}}, '{'{-25'd6486, -25'd3243, 25'd6486, 25'd1621, 25'd30806}, '{-25'd3243, 25'd4864, -25'd21078, -25'd24321, 25'd14592}, '{-25'd24321, -25'd11350, -25'd27564, -25'd11350, -25'd21078}, '{25'd6486, 25'd4864, -25'd9728, -25'd19457, -25'd12971}, '{25'd14592, -25'd11350, -25'd16214, -25'd9728, -25'd11350}}, '{'{25'd38913, 25'd30806, 25'd1621, 25'd29185, 25'd50263}, '{25'd21078, 25'd17835, 25'd9728, 25'd0, 25'd37292}, '{25'd34049, 25'd3243, 25'd1621, 25'd6486, 25'd25942}, '{25'd38913, 25'd16214, -25'd1621, 25'd1621, 25'd11350}, '{25'd29185, 25'd35671, -25'd1621, 25'd35671, 25'd32428}}, '{'{-25'd69720, -25'd71341, -25'd66477, -25'd51884, -25'd81069}, '{-25'd34049, -25'd45399, -25'd45399, -25'd56749, -25'd53506}, '{-25'd35671, -25'd38913, -25'd40535, -25'd25942, -25'd66477}, '{-25'd45399, -25'd34049, -25'd19457, -25'd43777, -25'd63234}, '{-25'd66477, -25'd58370, -25'd53506, -25'd66477, -25'd84312}}, '{'{25'd34049, 25'd9728, 25'd17835, 25'd29185, 25'd32428}, '{25'd17835, 25'd37292, 25'd4864, 25'd21078, 25'd9728}, '{25'd29185, 25'd27564, 25'd16214, 25'd1621, 25'd14592}, '{25'd11350, 25'd24321, 25'd21078, 25'd4864, 25'd12971}, '{-25'd6486, -25'd9728, -25'd3243, -25'd6486, -25'd1621}}, '{'{-25'd175110, -25'd145925, -25'd149168, -25'd144304, -25'd194567}, '{-25'd154032, -25'd118361, -25'd108633, -25'd123226, -25'd157275}, '{-25'd158896, -25'd119983, -25'd98905, -25'd102147, -25'd132954}, '{-25'd152411, -25'd111876, -25'd110254, -25'd124847, -25'd139439}, '{-25'd207538, -25'd154032, -25'd154032, -25'd145925, -25'd163760}}, '{'{25'd72962, 25'd40535, 25'd24321, 25'd16214, 25'd34049}, '{25'd34049, -25'd1621, -25'd4864, 25'd8107, 25'd9728}, '{25'd25942, -25'd3243, 25'd1621, 25'd1621, 25'd19457}, '{25'd17835, -25'd6486, -25'd8107, 25'd1621, 25'd19457}, '{25'd17835, 25'd19457, 25'd17835, 25'd9728, 25'd32428}}, '{'{25'd6486, 25'd19457, 25'd6486, -25'd6486, 25'd3243}, '{25'd11350, 25'd19457, -25'd6486, -25'd9728, 25'd19457}, '{25'd30806, 25'd3243, 25'd24321, 25'd9728, 25'd16214}, '{25'd0, 25'd11350, -25'd1621, 25'd3243, 25'd3243}, '{25'd25942, 25'd21078, 25'd4864, 25'd19457, 25'd4864}}, '{'{-25'd27564, -25'd37292, -25'd32428, -25'd43777, -25'd66477}, '{-25'd27564, -25'd29185, -25'd34049, -25'd24321, -25'd53506}, '{-25'd24321, -25'd42156, -25'd14592, -25'd43777, -25'd40535}, '{-25'd42156, -25'd40535, -25'd25942, -25'd32428, -25'd66477}, '{-25'd63234, -25'd53506, -25'd76205, -25'd76205, -25'd98905}}, '{'{-25'd19457, -25'd11350, -25'd22699, -25'd4864, -25'd24321}, '{-25'd8107, -25'd12971, 25'd8107, -25'd16214, -25'd11350}, '{-25'd6486, 25'd0, -25'd16214, -25'd14592, -25'd1621}, '{-25'd3243, -25'd17835, -25'd11350, -25'd16214, -25'd29185}, '{-25'd17835, -25'd1621, -25'd4864, -25'd24321, -25'd37292}}, '{'{-25'd71341, -25'd43777, -25'd43777, -25'd47020, -25'd37292}, '{-25'd71341, -25'd45399, -25'd25942, -25'd43777, -25'd48642}, '{-25'd71341, -25'd35671, -25'd22699, -25'd40535, -25'd34049}, '{-25'd45399, -25'd34049, -25'd22699, -25'd42156, -25'd48642}, '{-25'd22699, -25'd30806, -25'd16214, -25'd14592, -25'd9728}}, '{'{25'd29185, 25'd11350, 25'd9728, 25'd8107, 25'd14592}, '{25'd21078, 25'd11350, 25'd30806, 25'd12971, -25'd1621}, '{25'd12971, 25'd34049, 25'd19457, 25'd14592, 25'd6486}, '{25'd4864, 25'd19457, 25'd11350, 25'd9728, -25'd6486}, '{-25'd21078, -25'd16214, -25'd11350, 25'd1621, -25'd45399}}, '{'{-25'd89176, -25'd59991, -25'd47020, -25'd35671, -25'd79448}, '{-25'd71341, -25'd34049, -25'd22699, -25'd32428, -25'd43777}, '{-25'd53506, -25'd37292, -25'd29185, -25'd17835, -25'd37292}, '{-25'd55127, -25'd19457, -25'd29185, -25'd27564, -25'd63234}, '{-25'd84312, -25'd42156, -25'd43777, -25'd64856, -25'd79448}}, '{'{-25'd25942, -25'd29185, -25'd32428, -25'd34049, -25'd53506}, '{-25'd11350, -25'd24321, -25'd12971, -25'd22699, -25'd32428}, '{-25'd38913, -25'd22699, -25'd16214, -25'd16214, -25'd19457}, '{-25'd25942, -25'd9728, -25'd11350, -25'd22699, -25'd47020}, '{-25'd43777, -25'd14592, -25'd17835, -25'd22699, -25'd24321}}, '{'{-25'd134575, -25'd68098, -25'd50263, -25'd64856, -25'd118361}, '{-25'd81069, -25'd35671, -25'd19457, -25'd34049, -25'd82691}, '{-25'd69720, -25'd1621, -25'd1621, -25'd4864, -25'd68098}, '{-25'd85934, -25'd21078, -25'd27564, -25'd21078, -25'd87555}, '{-25'd137818, -25'd97283, -25'd77827, -25'd72962, -25'd129711}}, '{'{-25'd12971, 25'd8107, -25'd11350, 25'd6486, 25'd16214}, '{-25'd37292, -25'd12971, -25'd16214, 25'd1621, -25'd6486}, '{-25'd37292, -25'd1621, -25'd3243, 25'd6486, -25'd11350}, '{-25'd30806, -25'd8107, -25'd17835, -25'd21078, -25'd12971}, '{-25'd42156, -25'd16214, -25'd9728, -25'd19457, -25'd25942}}},
    '{'{'{-25'd147836, -25'd81968, -25'd81968, -25'd87823, -25'd127344}, '{-25'd102461, -25'd20492, -25'd38057, -25'd23420, -25'd81968}, '{-25'd115634, -25'd20492, -25'd21956, -25'd32202, -25'd100997}, '{-25'd105388, -25'd26347, -25'd48303, -25'd61476, -25'd93678}, '{-25'd169792, -25'd98069, -25'd83432, -25'd90751, -25'd152227}}, '{'{-25'd87823, -25'd30738, -25'd38057, -25'd45375, -25'd92215}, '{-25'd29274, -25'd2927, -25'd1464, 25'd0, -25'd77577}, '{-25'd52694, 25'd7319, 25'd10246, -25'd14637, -25'd76114}, '{-25'd52694, -25'd14637, -25'd13174, -25'd14637, -25'd83432}, '{-25'd112707, -25'd54158, -25'd39521, -25'd83432, -25'd161009}}, '{'{-25'd130271, -25'd103924, -25'd111243, -25'd64404, -25'd114170}, '{-25'd99533, -25'd64404, -25'd70259, -25'd39521, -25'd96606}, '{-25'd95142, -25'd100997, -25'd93678, -25'd62940, -25'd121489}, '{-25'd76114, -25'd84896, -25'd70259, -25'd58549, -25'd93678}, '{-25'd83432, -25'd81968, -25'd77577, -25'd55621, -25'd87823}}, '{'{-25'd24883, -25'd23420, -25'd42448, -25'd49767, -25'd127344}, '{-25'd10246, 25'd14637, 25'd13174, -25'd13174, -25'd55621}, '{25'd2927, 25'd8782, 25'd13174, 25'd2927, -25'd40984}, '{25'd4391, 25'd23420, 25'd8782, 25'd21956, -25'd39521}, '{-25'd8782, -25'd4391, -25'd17565, -25'd21956, -25'd70259}}, '{'{-25'd23420, -25'd20492, -25'd14637, -25'd36593, -25'd36593}, '{-25'd23420, -25'd10246, -25'd10246, -25'd23420, -25'd30738}, '{-25'd10246, -25'd13174, -25'd24883, -25'd2927, -25'd21956}, '{-25'd27811, -25'd2927, -25'd27811, -25'd17565, -25'd32202}, '{-25'd19028, -25'd26347, -25'd33666, -25'd23420, -25'd54158}}, '{'{-25'd80505, -25'd71722, -25'd57085, -25'd70259, -25'd92215}, '{-25'd58549, -25'd33666, -25'd33666, -25'd46839, -25'd65868}, '{-25'd35129, -25'd13174, -25'd26347, -25'd27811, -25'd60013}, '{-25'd52694, -25'd11710, -25'd17565, -25'd24883, -25'd62940}, '{-25'd71722, -25'd29274, -25'd38057, -25'd48303, -25'd67331}}, '{'{-25'd24883, -25'd19028, 25'd1464, -25'd20492, -25'd36593}, '{-25'd27811, -25'd5855, 25'd14637, -25'd7319, -25'd38057}, '{-25'd5855, -25'd4391, 25'd7319, 25'd16101, -25'd21956}, '{-25'd19028, -25'd10246, -25'd4391, 25'd0, -25'd42448}, '{-25'd52694, -25'd19028, -25'd36593, -25'd29274, -25'd67331}}, '{'{-25'd185893, -25'd134662, -25'd122953, -25'd108315, -25'd141981}, '{-25'd96606, -25'd71722, -25'd58549, -25'd57085, -25'd106852}, '{-25'd120025, -25'd62940, -25'd39521, -25'd61476, -25'd86360}, '{-25'd96606, -25'd68795, -25'd49767, -25'd58549, -25'd90751}, '{-25'd147836, -25'd109779, -25'd96606, -25'd79041, -25'd130271}}, '{'{-25'd60013, -25'd30738, -25'd19028, -25'd43912, -25'd70259}, '{-25'd57085, -25'd32202, -25'd19028, -25'd19028, -25'd43912}, '{-25'd64404, -25'd16101, -25'd13174, -25'd10246, -25'd61476}, '{-25'd81968, -25'd38057, -25'd27811, -25'd42448, -25'd67331}, '{-25'd87823, -25'd51230, -25'd60013, -25'd65868, -25'd86360}}, '{'{25'd48303, 25'd32202, 25'd13174, 25'd7319, 25'd14637}, '{25'd32202, 25'd11710, 25'd5855, 25'd23420, 25'd27811}, '{25'd5855, 25'd29274, -25'd10246, 25'd17565, 25'd16101}, '{-25'd4391, 25'd8782, 25'd0, 25'd8782, 25'd24883}, '{-25'd4391, 25'd16101, 25'd4391, -25'd1464, 25'd17565}}, '{'{-25'd11710, 25'd5855, 25'd30738, 25'd10246, -25'd8782}, '{25'd2927, 25'd39521, 25'd27811, 25'd40984, -25'd7319}, '{-25'd13174, 25'd26347, 25'd30738, 25'd16101, -25'd21956}, '{-25'd21956, 25'd17565, 25'd23420, 25'd33666, 25'd4391}, '{-25'd70259, -25'd13174, -25'd21956, -25'd36593, -25'd42448}}, '{'{-25'd117098, -25'd73186, -25'd71722, -25'd65868, -25'd103924}, '{-25'd58549, -25'd26347, -25'd8782, -25'd29274, -25'd54158}, '{-25'd49767, -25'd8782, -25'd2927, -25'd10246, -25'd49767}, '{-25'd57085, -25'd24883, 25'd10246, -25'd11710, -25'd51230}, '{-25'd86360, -25'd32202, -25'd30738, -25'd61476, -25'd76114}}, '{'{-25'd81968, -25'd46839, -25'd38057, -25'd45375, -25'd68795}, '{-25'd51230, -25'd20492, -25'd11710, -25'd8782, -25'd36593}, '{-25'd39521, 25'd8782, -25'd2927, -25'd14637, -25'd36593}, '{-25'd27811, 25'd4391, -25'd2927, -25'd26347, -25'd60013}, '{-25'd76114, -25'd61476, -25'd39521, -25'd48303, -25'd89287}}, '{'{25'd10246, 25'd5855, -25'd5855, 25'd4391, 25'd5855}, '{25'd1464, 25'd1464, 25'd5855, -25'd5855, -25'd5855}, '{-25'd8782, -25'd5855, -25'd16101, 25'd0, 25'd5855}, '{-25'd23420, -25'd20492, -25'd17565, -25'd20492, -25'd26347}, '{-25'd38057, -25'd45375, -25'd46839, -25'd49767, -25'd55621}}, '{'{25'd23420, 25'd23420, 25'd10246, 25'd4391, 25'd23420}, '{25'd19028, -25'd4391, -25'd16101, -25'd4391, 25'd10246}, '{-25'd10246, -25'd16101, -25'd19028, -25'd13174, 25'd7319}, '{-25'd1464, -25'd7319, -25'd19028, -25'd4391, 25'd8782}, '{-25'd16101, 25'd4391, -25'd26347, -25'd14637, -25'd11710}}, '{'{-25'd10246, -25'd7319, -25'd8782, -25'd23420, -25'd23420}, '{-25'd21956, -25'd16101, -25'd13174, -25'd27811, -25'd13174}, '{25'd1464, -25'd8782, -25'd11710, -25'd14637, -25'd23420}, '{-25'd26347, -25'd5855, -25'd27811, -25'd27811, -25'd35129}, '{-25'd40984, -25'd19028, -25'd21956, -25'd35129, -25'd30738}}, '{'{-25'd158082, -25'd105388, -25'd147836, -25'd133199, -25'd153691}, '{-25'd100997, -25'd55621, -25'd95142, -25'd80505, -25'd67331}, '{-25'd108315, -25'd89287, -25'd125880, -25'd90751, -25'd105388}, '{-25'd98069, -25'd83432, -25'd96606, -25'd77577, -25'd95142}, '{-25'd122953, -25'd89287, -25'd105388, -25'd102461, -25'd93678}}, '{'{25'd21956, 25'd30738, 25'd19028, 25'd80505, 25'd79041}, '{25'd42448, 25'd43912, 25'd21956, 25'd43912, 25'd61476}, '{25'd32202, 25'd27811, 25'd29274, 25'd48303, 25'd43912}, '{25'd45375, 25'd27811, 25'd36593, 25'd55621, 25'd42448}, '{25'd49767, 25'd42448, 25'd32202, 25'd43912, 25'd43912}}, '{'{25'd21956, 25'd29274, 25'd11710, 25'd27811, 25'd86360}, '{25'd55621, 25'd32202, 25'd21956, 25'd27811, 25'd58549}, '{25'd49767, 25'd13174, -25'd8782, 25'd10246, 25'd48303}, '{25'd42448, 25'd27811, 25'd2927, 25'd13174, 25'd48303}, '{25'd55621, 25'd40984, 25'd16101, 25'd30738, 25'd52694}}, '{'{-25'd67331, -25'd49767, -25'd35129, -25'd39521, -25'd70259}, '{-25'd60013, -25'd35129, -25'd13174, -25'd29274, -25'd45375}, '{-25'd51230, -25'd21956, -25'd32202, -25'd24883, -25'd39521}, '{-25'd65868, -25'd42448, -25'd16101, -25'd20492, -25'd61476}, '{-25'd68795, -25'd61476, -25'd35129, -25'd57085, -25'd74650}}, '{'{25'd38057, 25'd39521, 25'd46839, 25'd43912, 25'd62940}, '{25'd33666, 25'd38057, 25'd43912, 25'd32202, 25'd51230}, '{25'd35129, 25'd45375, 25'd36593, 25'd48303, 25'd55621}, '{25'd43912, 25'd45375, 25'd52694, 25'd54158, 25'd54158}, '{25'd67331, 25'd60013, 25'd48303, 25'd71722, 25'd70259}}, '{'{-25'd71722, -25'd55621, -25'd60013, -25'd40984, -25'd86360}, '{-25'd62940, -25'd19028, -25'd24883, -25'd10246, -25'd45375}, '{-25'd51230, -25'd24883, -25'd27811, -25'd8782, -25'd57085}, '{-25'd43912, -25'd32202, -25'd21956, -25'd20492, -25'd32202}, '{-25'd87823, -25'd36593, -25'd26347, -25'd23420, -25'd48303}}, '{'{25'd45375, 25'd52694, 25'd38057, 25'd24883, 25'd40984}, '{25'd20492, 25'd38057, 25'd27811, 25'd13174, 25'd35129}, '{25'd14637, 25'd7319, 25'd16101, 25'd5855, 25'd23420}, '{-25'd1464, -25'd5855, 25'd11710, -25'd4391, 25'd38057}, '{-25'd17565, -25'd27811, -25'd24883, -25'd8782, 25'd4391}}, '{'{-25'd61476, -25'd45375, -25'd54158, -25'd64404, -25'd111243}, '{-25'd13174, 25'd10246, 25'd16101, -25'd1464, -25'd52694}, '{-25'd21956, 25'd5855, -25'd2927, -25'd14637, -25'd48303}, '{-25'd36593, 25'd2927, 25'd5855, -25'd17565, -25'd46839}, '{-25'd35129, -25'd35129, -25'd35129, -25'd42448, -25'd79041}}, '{'{-25'd14637, 25'd0, -25'd19028, -25'd32202, -25'd71722}, '{-25'd17565, 25'd14637, -25'd2927, -25'd14637, -25'd51230}, '{25'd0, 25'd2927, 25'd14637, -25'd1464, -25'd43912}, '{-25'd7319, -25'd2927, 25'd11710, 25'd4391, -25'd49767}, '{-25'd26347, -25'd20492, -25'd29274, -25'd21956, -25'd65868}}, '{'{-25'd36593, -25'd11710, -25'd23420, -25'd14637, -25'd27811}, '{-25'd10246, -25'd23420, -25'd8782, -25'd11710, -25'd16101}, '{-25'd4391, -25'd24883, -25'd4391, -25'd5855, -25'd11710}, '{-25'd36593, -25'd5855, -25'd26347, -25'd21956, -25'd39521}, '{-25'd29274, -25'd11710, -25'd19028, -25'd23420, -25'd32202}}, '{'{-25'd51230, -25'd23420, -25'd24883, -25'd13174, -25'd30738}, '{-25'd23420, -25'd10246, -25'd14637, -25'd27811, -25'd17565}, '{-25'd38057, -25'd23420, -25'd30738, -25'd20492, -25'd45375}, '{-25'd27811, -25'd10246, -25'd20492, -25'd14637, -25'd19028}, '{-25'd19028, 25'd2927, 25'd5855, 25'd11710, 25'd4391}}, '{'{-25'd51230, -25'd20492, -25'd32202, -25'd27811, -25'd65868}, '{-25'd38057, 25'd8782, 25'd2927, 25'd7319, -25'd29274}, '{-25'd26347, -25'd4391, -25'd10246, -25'd2927, -25'd51230}, '{-25'd29274, -25'd1464, 25'd4391, -25'd29274, -25'd57085}, '{-25'd84896, -25'd58549, -25'd55621, -25'd43912, -25'd79041}}, '{'{-25'd67331, -25'd55621, -25'd20492, -25'd52694, -25'd62940}, '{-25'd54158, -25'd35129, -25'd16101, -25'd17565, -25'd45375}, '{-25'd38057, -25'd16101, -25'd11710, -25'd13174, -25'd40984}, '{-25'd62940, -25'd29274, -25'd19028, -25'd30738, -25'd49767}, '{-25'd79041, -25'd46839, -25'd39521, -25'd43912, -25'd74650}}, '{'{25'd5855, 25'd11710, -25'd13174, 25'd11710, -25'd10246}, '{25'd2927, 25'd0, 25'd8782, -25'd8782, -25'd24883}, '{-25'd1464, -25'd8782, 25'd16101, 25'd7319, -25'd19028}, '{-25'd7319, 25'd1464, 25'd10246, -25'd5855, -25'd13174}, '{-25'd11710, -25'd11710, -25'd4391, -25'd16101, -25'd17565}}, '{'{-25'd65868, -25'd33666, -25'd36593, -25'd60013, -25'd95142}, '{-25'd29274, -25'd11710, -25'd2927, -25'd32202, -25'd46839}, '{-25'd7319, -25'd1464, 25'd21956, 25'd11710, -25'd32202}, '{-25'd24883, 25'd1464, 25'd5855, -25'd17565, -25'd49767}, '{-25'd51230, -25'd14637, -25'd13174, -25'd33666, -25'd58549}}, '{'{-25'd98069, -25'd45375, -25'd38057, -25'd62940, -25'd62940}, '{-25'd65868, -25'd13174, -25'd2927, -25'd16101, -25'd45375}, '{-25'd57085, -25'd1464, -25'd20492, -25'd23420, -25'd49767}, '{-25'd60013, 25'd5855, -25'd5855, -25'd33666, -25'd42448}, '{-25'd89287, -25'd51230, -25'd27811, -25'd65868, -25'd92215}}}
};
